-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
T+H7dX465QawZm03xg+n4JsPd9TYeUVmN22UF96eoBBqImseipOMK4YGsVLtcve1eQNTn+oWjVnD
9UZMKxPxf77mQsNSuJ7hj0q9uPH0MMLZ9pd34r8wGDs5+d0Wkyklv7j+66la6guqrvYThJdy0ir2
SfyeQiKOoDxEdfZ7VDF97gaRFyfLL2m3TmER9TxmH3TUq3B8GvayHPQXpE22IDUnTWaOZkK3q+Um
kvhQqaS1VXZNGJFht7J6VEB6ZFvVNJwN0RAPvSmMnbK0FbAFNngbbVhW1dvIZONe49QwKjXuB/t7
Xy+iOGhEjXK3vTVCK+S9oPesZtxD6+qSsFO0Kw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 1072)
`protect data_block
ssAoVO/X4Ov9AeRz9Kk2VOgD8V5u1j9tlDsnpTkPeCn3EApiVr5THWMaQ2EBgyfMpXJqiVCVf8BH
qiDU7wd5+5yGX8IDzZLcBrcpNsSmH3EtuGc071zxs5J/v+Ws4s4XZ/VLqCwwfbrIW+bKYAZzKk/D
cow1IFcYeiP3OBAwRI1iZo14k9tPNe7GGhz1fAz4Pi44uDo6h33tGSBNBdnwFOwGCBz85r2Rll7p
r2WNMtYbpJ8ZsrhjxzqSU1S9XAa9vxH7G1LuPcxzzDM4Z6044w/onfOCvcmGmmGbhGmt7JxOJ5KR
xuIZtUfszjdlU0uWp5lgY7fW3w0ZGBhbH7Nz40O4gaFRzu8iu4VciN6kVcWr2IpZeI2t/OydhfsH
q6KyhBxrZVx+21DDHSx5AVqZ9I8ekr9yfScDRYxNV8G+xPfcmWq9mgd3SGhjYCoTCnqZ/sqgklwx
oSL3/UpHJgubhUxCji3pdKUzsyFI6PpZls8wNbQo2RW7h4kBeqWDKRzBNCWPRgSH60XwmXiRR7E/
xnouyx9HaA1nFGv/2xmBpCVPwkWR6n1RsHbvHJi+oMhKgOinkQGJEtpFTLYN8QmAxwom9Ewu2uQq
LKUOFnSGKADl8H6i8X4+sxRTK6EcovCDGzQv9dQJYKctvv/+JwO5squerP/CjiewOIJ+YpVAq0pC
mflHfxLgep131ZeHrWUZr16gFSSqwKW7e/LRvyj/DqCB08+6s4pWaEfXzN8vEuy0a9M2ce+cKGKg
7j8w39RalMVmgpfDmHSWVvdgdnzrlLV08Uyu13iwVOmLnfwo+pwvqoGlyOYqZA+Ex3R/Srm01j4f
J3Ozcv2uYBIPyql0+KvwCf6MvQZEVGAuPAWQ+7tjcwMaM4DB6R3KX++zQTVpK0+GVRB8JQsSdTqK
W7VWjb8eF4qWkbFh8/T4IicNoyQQnOawN6TryvssoLBBpFqHLyLu2VaSioS2Gk71cVLZjuaFsTmh
aGEUwtKLGI2+sskdh2RLiRkAkBaol8tCcz0hXQdw8B9X4q1/TzaWFTQa/oRjbyQI9+3SXPk6uZVn
kH/sMZeMXAkJ5O+1sOtrIkTszP2ib+6376dc/+NlFoGzlAWhPJLA/gKQs0mdhnuHW7q/YgzFqHv6
IQsd4zQP+Torm7glusNSkMfwLZzGfUqQAZ7xt3PhV5l20eNvO6XGMlSe8lXzTo8f/zEDipoHjjl9
37C5VXXMWfPwWDmryepA/aoQhXRXN3hNe/TuCOdQpXwRzUm45FBgiC2+s5840ELEnOubsMUL77Av
reozh757y3XEo0B7aracYBglY8RLQAn5PDMUcX1qet441Llm+XUMUnkdCbgUMLYj7EtbXm5aNGIn
uQCuURreoQyoQN9zWBDS7wiWecUqaf58/iXYQpdSzeCr0kKFdnhuKJxDKSVlfw==
`protect end_protected
