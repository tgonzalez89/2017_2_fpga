��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,�Q����ф�74$~�I#���q=6�;rN�/O��<�qAC$,C����]�-���^�o��5,A�X���5g��|���Y��z��� q@�[I������C9��"���c @�W�-�8�����փ��'~����VX���#�)p�>�O52==�SL'?�u��L��׳b����~����w@�"�ˏ�IW��'[�j����`����5�Z8�Xǿz/��
\�q ��P��7�B��䌮��a�Z؊�S��Y�-+���j��\=)�[��2���K�g���og~��2��ן���lP�ad�ĊT��0$_/��|t*�e������m��7H�Y�)�LQ�u�m��|��~p��+i�}(³ߣ�bJ�3�\�����٦l+g�X���ݘl�_$g�_~p�8]M8le5SiL�r�vҔ����_9��X6md��'=������ t&�_=�h"����H��8������j��V<�N�.r)o� Y�[��-��������) e�%�S��W!We�g��1�Ч��\��!� U�
��(������_����L7XS�?@'j�"B�h��� ��mtmSӘF�Z?YXp)d[ڪ�����t�%�}��<r�ѓ@�b	�A��<1\���kiq���Cy��;ِGy0�wz!�Z��B��кe��.�a60)��@�pɀ�&3G-�v��~Mij�����W�6�X��^"&2Xa���X���Cɴ��R+�ꩱ�!RU��z(��:֎�:�}�0�p j���n�E��Pe�~��m޵�Cn�t@�|@�ݤ}����Mc��y=]��j�{�Uհ�.;��8��n���o�j�|��dh$2�0J��%8q1A1$��Xf5�^�z���Gxl�Y֬���k�]�4����K�d=? 8yҦ�6��r�<��pO[  �	m��QO�&�e�x!X#|�j�����'�V� Ҿkhk�).�	K�{�A*]Fx�S�[��,`�H�+�W������`Zx�-�vX��n��ں� A���������.'�}����ϙ����G��ϡ����͸`���VX3��&��4>�q��$UYQ,�1����X͋52��3𐒈e�{�+)��
�y+�S!**�<7��q�T3�s��2&��]~-;�0�����>�6�B��9���󼃒�%� ���s�Q�2w���J����l�C8�'��L���_T�L��yk��W"�/N��uJB�]e(���y�x����7�h��|����d�-�j�D��a���YƷ���G���#�nH L�������(H�����(:�d����_��f��^��F���G�Oz�MZR��BUm������kr�l�W�a����m�ʭ�yp�)�,���`+�R�o��Zg��84��3�A�S9C~�C�mMp[3(��u��p�)y8����wD�n5����q�������榞�%�Ik*��Q��`�	P^�r2�h||=�~����O�	Q�Hh���=Iuޖ*�=�XCi�ɗ�D�D�c��� h��F�b�w�̊�J�%|�7�5���Daub�O�/֩�$� K~d�^qU2͑�iYɽ�e�X�$gY5�b� )��K�d��z��+Mm˖����dm��Z�s�8��t�o�)p� ���2�9��H�y&o��rz/���~sW��_�ǐ./+,i���e���,q3�`t;X��/?#��e���/y���#�Z���w�uɧ>�D�(�'�oV	��+��z�p���y �wU��H��q%�*�S�BB�H���R>^=7��$�5�m�3�kdl�2˱�2��d�A?���I�%�3x0.�V��o7����2���ĉ{�u��F�K��"��4�ż�~�\G�{(�b�a��!g&��4�̰�j�zz�����ZD4U�VF��l�E>���f�W^)`9�{pQ!I��b��$|<\�.{�4᪱���U������#�8cZY��K�g=���@y��6����A�.��C`�T��ǆ�v��`�L�n���֘�=4�wvn$t���r���P�GJ�����>�R6�P������@�����r���B�J�[��B��#������|u����3����Q��Ej\(����8#��j,�t�lOo�g�����	Խ:'XҍSU|t�X�.�.=�.}�:	�%V�ea`�����0��"�q !l�˩��e�G|�|\0�D�"�U��"Pj�N2���'���[O���/�{À:��U�Bs���d��5vqXa1�}`�{�ZRD�3��/�2sc��v�VzBq��."L��T*G_� � �C^Pذ�a� �_e	��M��s��M�������r+2C�]kvt��R��$t�v^`n��n[�6�B$٤�:�!bיF���y�K)Y`���´K8�
��x��/m�R���
�]ԡ���h`�q�L~0�Y����e��Ŧ����b��
�oɷs*�a7�q�Tb�fH��sf���O�G�C�kO!����˳��M�^��&�%�B��K1��b7�qaC�Zf�o��O#o�0^�DV��i9Wa����"�ђS)���1������y>}�<��X�|��!C|d�25�9Miᇏ8��!��*��W��6��3 �7uA%�-�XS��