// Copyright (C) 2017  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Intel and sold by Intel or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// Generated by Quartus Prime Version 16.1.2 Build 203 01/18/2017 SJ Lite Edition
// Created on Wed Jun 21 17:54:30 2017

// synthesis message_off 10175

`timescale 1ns/1ns

module FSM_gen (
    clock,reset,tx_almost_full,
    data_sel,tx_load,fifo_rx_read_rq,CS);

    input clock;
    input reset;
    input tx_almost_full;
    tri0 reset;
    tri0 tx_almost_full;
    output data_sel;
    output tx_load;
    output fifo_rx_read_rq;
    output CS;
    reg data_sel;
    reg tx_load;
    reg fifo_rx_read_rq;
    reg CS;
    reg [3:0] fstate;
    reg [3:0] reg_fstate;
    parameter IDLE=0,A=1,B=2,C=3;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or tx_almost_full)
    begin
        if (reset) begin
            reg_fstate <= IDLE;
            data_sel <= 1'b0;
            tx_load <= 1'b0;
            fifo_rx_read_rq <= 1'b0;
            CS <= 1'b0;
        end
        else begin
            data_sel <= 1'b0;
            tx_load <= 1'b0;
            fifo_rx_read_rq <= 1'b0;
            CS <= 1'b0;
            case (fstate)
                IDLE: begin
                    if ((tx_almost_full == 1'b0))
                        reg_fstate <= IDLE;
                    else if ((tx_almost_full == 1'b1))
                        reg_fstate <= A;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= IDLE;

                    CS <= 1'b1;

                    fifo_rx_read_rq <= 1'b0;

                    tx_load <= 1'b1;

                    data_sel <= 1'b0;
                end
                A: begin
                    reg_fstate <= B;

                    CS <= 1'b0;

                    fifo_rx_read_rq <= 1'b0;

                    tx_load <= 1'b0;

                    data_sel <= 1'b0;
                end
                B: begin
                    reg_fstate <= C;

                    CS <= 1'b0;

                    fifo_rx_read_rq <= 1'b0;

                    tx_load <= 1'b1;

                    data_sel <= 1'b0;
                end
                C: begin
                    reg_fstate <= IDLE;

                    CS <= 1'b0;

                    fifo_rx_read_rq <= 1'b1;

                    tx_load <= 1'b0;

                    data_sel <= 1'b0;
                end
                default: begin
                    data_sel <= 1'bx;
                    tx_load <= 1'bx;
                    fifo_rx_read_rq <= 1'bx;
                    CS <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // FSM_gen
