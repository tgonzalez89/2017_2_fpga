��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR���[{�T���CK��TC,���:�
&��d!��]9�'D`�"9 S%�aQ�`!�6������V�W�l�a锦E(�\gC�slu�4U5=1�N�m��l�9ў��P���B�@+yg��=�}|֦���ָJ�,������
���NPx�x��b�dD��O�+3� �	�a�?���9��b��?y~XW^D\�>��GJ;�ߏ/��׭����wD�%1�z-�Ϫ]�޼6΅����Ĺ�}��@�D�O��CO�$�m;y]�x��!�}��~���)����RQ�0����£5�%��xV�"����-�{���],FX�^�>�oh�}zY)M�T�ކRk��z��%�Ep*A#�}��c'ɂ�1�B҂� @/tJJ�
�K���#���i,E՚v�Zq���géԃ��9)�E�!_$JKj\�,F�X|�]yt**�K������#�2�?^7}��%��b��)��=��Z;��%���'Nw~���l;�;||2�l��Ws�	d�+y�(�����Δ�ZP�$�ܭf����Nh�����H��h,�N`��{ڏ�O��L�� 6Ũg�����\��1�?� /���f|v���v?�Y�nw��}�@Saʣ?蘟�K(���׆���D�r��+��,l4����N2b�?�$��#%R���Z}�Jvu�Z�9��&2EZH�3���El*fX���ճ�Y��dk\y:��g9Wlu�*��dZ(�"&�W�|JeS�i��X����%=�����G�<υ��ǭ��6�\L�M�1�Qs)���ۈqƄ��޸��[�D�0�e6����`oc�D��S̰%�𥀥�*Uw�,����jDHW8�\�u�8ݳb��ɰP[�����T��6��W3�T
�"t5��~AI�����<�޳V!=��y�ŭ�k�DB!u������g��e7�����g0}㝁��F��[AU���oQ|��U:(�
%Ty=g66��"���Ѽ�I��ˁ\��U+� ��fH�����X6e�Ɋj@M��w��Se�At�3o�ݠ5�U��!���M���,M$7���!MB���\~")���������2�)�Ȟ�ȴ Ǩ�&g;�DM��"rwB�5��}�Ճ��536_iѣ���r���xTg>X���"8م�u�ܐ��i��2��)3+�s����%): Nt;$#���~�:��W��`�`,�!�.w�*��_t?����Od�Ū!O�3�z�|�O�g����·������Ֆa��f��{��i�e���T�|MT���f˭����z7�כT��LFﲇ������G,�[6W �j�=�@�|��c�Q_���$�x�ڰ�GKɾ�>s���s��bgh4paqB3Qwјz��^��4�l�����י�n��e:���3�Fe��$u�2���,u/�6�2��9c���[>`AŀpFk�qe�ⴐ�F�6�0�ȠM�&�٦c*aONT�8Q��.$�"Q��5�R�Pi'$��3H��:�xg�	�6�R��5����V/�7�@�=�OY")pp�c�ρ�n+�pWt&�m�J�혈�J����7t.��bV"@X�Ե)�ߐ���m�s)KS���
�s5���e�#	1��'`.<&�:B�wgM�#p�q� .Dz<Mx��v�C�8.�;��o_�>�3{Z���,���]��
��۪ԟ��{�@��%�7.������]˥��v�W�w��k���P�6���PXEj�>�[_z������	�#��������!T�#}A��&�3{�h�?�v	���y+�_�қP��l��M.P��N� �)/ꗻ!���)+��h�]ۋ�L��d�{K�\r��s0�
H�_��B�:c��~�b�?��_�s<IU�4�KZ��+���L��~f��L���s�5u�z�s�>ތ`���V��ʯUOk}cp1Ίq�X)�'�j]�қ�������C�(�L\RY��s�O�ۈ	c�� �{���4�z��;Iy��4"6��r[��w����U�m}�I��2�h�ӳ���!�����lC������~bG��U�5-54Ґ��Gh��Zs�i�TA�<�ш AX�K�����oYPl�O��yq��>���zd��oo{9���y��[�q�Y�m��'!��v�Bo%)ܨ݊��hIm���d���;�-�A �N���'3�v��=�Aߕ�+R��˸y�gp���L�6�{8�x���L�낲�6H�lH�����]ʅ��~y��H�T
3c	��-&�i,{o���&�+�dqm�͗����y=y��cZ����*B�-�л<�C��
;'��B��#���Z�H���P�ڲ�pWť0A�)s��F����0]���3I6�2#��A8a�oܻm8� ��/�RJ?�"��Ft��]ĚFN%N	a���[ի|�d�f�閞���[,��\`���kH�R\2lf�u��H������I3�uC/�G>�l�a�&�JMA*�+���C�?�⹠����+���*5���'/2_/�AL�Sv[���G����e�������Y!0��ׅ�-��J!��d<�$$�׫��C��6��[wM:��:�Br�����9�C64R����$��/P�_��9�Ӫb+6�@n�z4"��G��-��Nq}/ҀC����T��'����� ��7�㒀e����qh�j������٦�c�QP�[�v��a=��J@>�Z���T?#�xy7��.�#�9�<j�X���� #8���}Q���O��C���y�g<FBJ�wx�G�zʒ�?��3wH� ��������)!C�/�U�έ�d��_A�t�~�C�ߜ��x.�?WK��N��e=*��{�B+�B�W�bO�^P:p���	��W���cuve+�T�����/�;����J�W4Wjf��*J<���0,�hH��)y���cX�#�SP�X���,�̺9��)���)}�a��/3fN��yp�{^�����j�f|��
%
z��H�N7g�d\p��0���/5*$ I
�'n�k�<�Az���H�p����%T�=&�������T:F�O,y��C��v%i�P�ɜJ��.��U��A�����X��:�%��?�\e�1h�2_x����������~]��N^2S=Ox����������-됽J�y���v�1��(6�olg�[��!)2?`l��ٌ\]�;a2mw���=��(��jHݴ�����t��o�L�돘Q�����3��Jb��-�N�	�I����*�����[���m��Τ�_K�h0Y�T>��#��:�Of�����������$Շ�h��G�Z�+�ӡD�R�%=0#�T:Ŕ+~S�q�����b��u�N��?\���T���Gu������,��R��aR"9b�`��Hxt\L�F)�
&�qs�b5��x76���i*M��&"�e���x���k�_��[
6�������A��|1�����o��-�ɦsfc