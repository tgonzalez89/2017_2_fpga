��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,�Ȅ���P�#�J���zzJ3~,M&�pE� s���sH6�s#>_y�}�j�q�j�2:K*��j�,��
܌r���ҷ����&��)U�����f�4��	s����9	� �� 2)��.�'�����^t=��NW>��xU%�*«e���k��*uvXN��z=6���=L��ɝS�~�v|Pm�Z��0SOc���}&;�gu��cy8�f�K:n���pP��	�n���>y�)���h����И?5���Zdu��ީ.�2wE�C(@�+!~*o�	�� Ԛ������2��acg�����B�gI��5��;�p�� �1����F��߶f4>�y��&�K^n��WD��'���kA���`����b��s�]�_�TY\@F]��̸]�V2ު�܃��&
"�G�Rb#l���C�b[�s��� �&��.
7e��o.QmHx�e^����r���
˄�ݵ���C���!FC����"Y�#�ٗ�=nO.]��sW~��J�iGV��'�����KR֔kP"�+T9ݻGR%ɂ\UC�'��k6iԦηxp��$9	�=r�"v;5,�E w�%�H�Sm�I:8�W�S! ����]�����O�t	�zF�%�1+�d�c<w�0sJ���/*s4��n����30*�ᑽ�J���x_�N�,Wi��t,Gz��Ƽ���sⴰ�i��������w�@x�]�&�%E;��%|��qOHu���4!�Q?\���� �,쇀�3�MAF[	Xx}3/N�bP���^l�Y���^%�~f���^�Ǚ�4�,bk[{y{�d]�斃���0}m�[I�!jWO�ޭ� �eAo�s�7Y�4��E������$3�e5aU��u0vJ0!��(�Q{�������3M� 7�����VI�����f+��?ܶ�㔀C�5A�0��-�$q�Q�(*���-wm�r�Tc����\�hy,Q�i|���9Hl���g$�F�4Ms�w�� 6�C/�"J���$��73}�����9����<�!(ʞH�'�u�wB&A�4��)ن�f��3|5�ta�xx��Z��h\��<dTA'Cr
�3"w<-풼"��*M�Ȧ�,��H|<�}u��D��b"$��Y~t8mxD\O��8�J�����/�AS�:#�R�zg(��4K�������J��.,^g��p��fI��;-Śn(W��(�U�]��E�|��*��p�;�;���S�G��%R���y�
n�fT��rH�?�䘺�R�v�{�l�����{�M�:�X����`��\���C���f��u�oU�J�n�D� y���|8��j�7�<� �#�7������b��ǎވ8R���\Wu4"��86�j������;�F�4��r\#����q��Vmb�m�"��9���}O.R����*GSO�K��S�֠=T
u%�q@�w�6(�`[����C�զ�n䶑5|���w��x�3��w|j��o^�$�M3u*.AN�B԰O4&�eޒ����RK����yTU������+.��t�ʳ��0�/��o��i]�������(ƫ^b�7��gD��f xP�j�S;c�j�ӯ����3���J��W��3�sFk��=\�"s2�,�bǸ"��Ȣ0�ϗ�(�)��}���SwY&ss�_ܷ�(톳� �\�1�u|��"�7?P/y����8~�٣��Yz~b+�Z�X���Ys�!�V�!j�a8��oB���꯫^F����u6�3����黱�����4���r}|�&l'�8,�t�;�5��PHZF�6.�{����3n֙0�e�m�$��{��P�!��޲�M��caʞ�&�N��w0hf`*�C!�S��W�O��p#��I�p��A8֟�߈�C6�'��Lm�x�K�4��Eu���1VH
)���x�z�&M��S1}��(1zTlr�z�
�&ގLIdLyCM�d���|vr?]�3���K�y�]XfC;*S�uͤѣ���0j��vGI�d�R���0t��fj����w��~��_��f�ѫQf�]�>1+�0�"�a.�ץ��&�aȕ�hk'���|�_ �0�ai \������H��v��¾�z%��E���u�B�����ㄗU@S�C�hͶٽE��tS��C�&��!�㢃�%7ܣx��(D�oBx�.(Z�hT,��✦��X2b}�kh3��b�7�-}�� �Z/V�4��L�
!.=13��~�`";l��7�}���G_�'G���s��E�~|�[3�-���L�~פl�����d�t���� -ѣ(Ϸt7�S�Տ������Nl����������9��K�[|�� :xJ���v�U8�ƽ�;�/�G?ji�
��u�6�F8г��w�]�(��pŮ+��%�Õ�ο���D�n���h.`�HQ^>���/�M������Ķ��	�5���3pXӹ}�����~�\�c��	�@"��$5��X�C^���+����FH�kW%��5WG������xԸ�ġi,��i�Q��B�M�O��j`�)ӫ2�� z��#]PO�d_�z��U��FP��b��=�.�W�r/2���L9S��L����͔�fr����O��z#~1@N�	��
FL�~xو�!���|#��jA�Ob�ܽ*��p �n7�H=�L��_%�P�^-|��qa��oˑ�7A�T����g�&�W�Y��nd��WҮ0i�ڹ�-%��������d��l��~W��0Oo�}��7U�Rڶ��9��F+i��)�#	����1-�a��,!�p�/f|�@.kY��6���ǯH���a����+�{c.T�tW7�Y���n�Yϫ��,c��#�O�}��1��|���z�?y߲��1�C�I��p2<�w�u��I�-�mc�Bx��)O8��#<Y;r�27Ͱ�{Y�d7�*��UF�S�D�?P���L���Yl�s�@�
��J���%c�����\*2��}[:Sܝ��G
-�J-U+K>|�$f�;T�}&цm��kޤO��8��IU����Hs`�-���î2�P�-%�d ���ʍ�M�l�CeA�]aL��R�����$`a*X�u�f��X�W��لШ�Ú��w.�8� ��amn %��E��f���M����aV0&A�8@m"����Vdk�8��3�D��6����Ϭd����v�F\��(��~P�ڦ����G[���u�1x��������tL
t�ۚ�H�X��mm����Tw���ƪ�w�Z��+��2�A+�οaZl�0�A�B{<?꒔�?h�������������e�U�h��FLU\��/��{��Ÿ�Pz 2���DWЁG?ۨ�d	��-�ܰ�ՍU�$��`�^����QJ�eq���8��6�9y�^j'�+�����l��4�!N�hC�Zב\���F>���c�s�$��B�Y6Uj��ObQ>��3� �g+O��
A9��q� �A�e6���(�R�r�ˢ����[_�,�����k�̝�ݴ���Cv�a�p�FiW��w@����K��\Y Gw\s9)�n|�ao���x��4ZL�t�׏<�mO�a&z�8��~4v�ZH�G����+�A@�bwHq�\���-�&6�y��4~�=6�aNW��,�>�d�˰�'�mP���5=���@�������Z��mNҌ{�"���&� �D���qT��X���)����%x�F��P�7�ڿ�01�f=ΖǙ9�I��	�p�i.��GǑ	�d���i��VYH6�:8p��r�t\K���|X��qg��تu��BY9�V��#���=���� �vt�f�OE�M���D���n F|��bC��-u/�D#t�"�P ��
=��u6�{M���	 А�G���X����e���ز�3W��yY�Բ=p,6{`.��&������zP<(	���;}�ޥD�����͙��'��8�}Ȅ�V!�R�r���jf����+8f�ۖ��m�ɲ�O����<x!]7�)�e=�� ]�:J�Y�^��5�2I#%pq���fq��h�W�U��]�82�e3n~t�)9�m�2�@�igԔ��E����Q��#�R�P�<�ʁ�ͼ":�S�����<	�g��THX��N ;,�>|�}�<��Pf!=93�:1��Y`+ӕ�/�I�ޟ��;`}=���k̈��Ҥ�D��,޴!�ȑ���N�N�����̿�^&��n�쇪��7:#���)�P����co���PD����/z��l�H�u�Z���lJ�$�����������s|Y�h������׳h����e=�i�;�d�4�2�@J�u��5紨ć{����t�pB*B���H�T��!�_M=i7��o�|jC�f#�d�j��Q#h�Z>��)�|�5�t�J$XG��b�]�>q
�����x� 2aY�eͶ�E��tt��,��Q>�i~�xa7V�e	��"��#f o��6f�4<!�k,Dr�P9� �C-��}�����V4㐟��Ō$��]5�F*�,�`��V%��3,Ы�̌��G�����7��C��;��/}>CN��wkhE,�) ȓt?Rwɰ��jda�(Goܿc25r/�|�_�+�U�۶5�ө)-P�rN���dec�h�W�Ҡ���&�BvI���[Uc���uH�o��X�f2@FeYlx-jys,$Α�/W���ŕf�7�+M򢄤{�x个�2�P�_���9����-"����*��"�S�*L���>V����ʸ�K|�ִ��^xd�Hzj#U��\~�,�PR"h�Ԑ�z�HJ����.<�nCC��L��YQ�[ƭ��nH�$�S`>
�x�%���b���|`޵k�̜K���^��J
Dkou�Y���-��jjS/2�X�O� ������E#�~��iY���}��>���z��W.7C5�@<&�(����Y�J_�2mP�%��N��-�=��c�l��HOS��᧚�F�W]HO��M8X�x��
�zZ�(���,Mq��¦fm�U�/�!zPJŕYL~cYL�!�k5Z$���j?^�_�'���t�t����G��}ִ�,z�� -���KX�y�Fb�oQ⤛�(`�v�"�1�y�̳�����f�"���Y�>E}�)�r�|lh�<���Mh����+��ٜ~b�c�,��u]�3:�9V��DW�7����4s����]p�!X_1�G�g�ix�R��u7�ңv��-ܒ7���[pOBO�(YҸ�S*qh9�8���������7ck	��w9~�)S����`��=� �q��D��Q���S(/b�s�a �Y�s�X�����J��DiW�����[��`ϑ¦c�]@n��r��<�VW��(rQ�&�P�>l�9�Y�9Q�:�B�Y���PqD��*�%~=�n�\s���h�7&J��[d�D1��%���'k׫����I�?�@���t����cQ�'��"1H*�ҴII�O���Su�b�`'�[