��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR���[{�T���CK��TC,���:�
&��d!��]9�'D`�"9 S%�aQ�`!�6������V�W�l�a锦E(�\gC�slu�4U5=1�N�m��l�9ў��P���B�@+yg��=�}|֦���ָJ ���;Qx�Y��JN�D��ֆ��@�� ]P���a�QYd�w [pى�[�{��B�y�-4@3m�-��Go�f���=��%=
�����	�M�OEZ����$HE��X=o�����ʛ��~5���|��q"����wG0b?M;*��� ����|�w����� ���>$9L��Ѱ{%_-���p3�\� ���|�J�o~�i�x��6�R��Ӟ%g�+\"v f:�>85+�ojs�eu�[��>��Vq���@���D7b�,IA�a�S��G�\��F\8$������m^3�dAe���i�tW�?��b3����
C-���'���UX�3G�;�e�(\���:���<K7��mN���bL����� t<u�tF�&�S��O<ǰ��a�A�R�9d��1j�4���R(�`�3h��g�c�{���J�Y�(�/�`A�)j"W��4#Ŀ	˛^H���1���d9�z-�F�'���VE(��4�o����l�>�ܫ���
.��ѸP��`c�������n @4H�8��=�켖��M� C���]��������n������2��|��x. �v����5�7�QĿ� �sq���;�&z>��4����s��~��3Y�I�Y�t��c��Uw@�c��a��^�����N����Ǣ�,z�j�|YOS]O����\�	U������
�S��#�@z��.X{�f�G$��p^#%((�	[������9�.�Db���.g��*��l����WI�.�r�ĪC��hQq|����
 XƄ=(��}�¸V�V���V3}ʠ���T���*-��uY��&��s�F���-��i��gQY\HH&��g'��Ms��d�KHlڿ���*�;�m�2���#5"S�l���8띕I#S`$MًQ۴I��P��1#j $��Wq*Jk�F��,��'6{ٍz�W I����B!z�8V�"�v�����u_O�����!���Aԫ~����h�T,�
��Tf�?��|`�2��!TGIL�]->��" !gUsF��v)�Z4R� �I�� ��(��ڵ�̍K��q; }�%Jzꆑ�?�ŝ��z�O��݋L}g��}C�j@]��!��������dKY���479O`���5c.��6��6
��+�ӠD���.`����L����B��w;��H)g��u��7:�*9�����E� R��㇘��}�_u�xך�*���z���	�"H�#.�<j+#�ot�M�ZW�F��ڵq�K@|Y��ژ m�?81P�/�=z���ɲ�X4MQKq�K�����;"�"�O
8��gH0͑+N
ju�����2�Ί���Y�Y�t#�R�Em4��[%��L(;+���� ��@�F=�r��Z'� �2�|��9�:Mp�f��<�΋���ɜ�$�=<�p��&U_wC�9m�ztcw^�)p�J��J�o�[�Q`񴴇<C�T$�_}�&I�٭1_�.�a�%h'2��W�zLʛŅm�tؿ�#�СA��@w(��u��4�2���]�'�d�>��դ�7�6�Ɨ��|��˛mSHʸ�GL�
=��X6.{v��h�I�������q���-�ד�'/R�-��u?����$�2)́8q�G`�0�!�0���R�G���Hɦq#y�(��t��.톥��ז�'�i+���|��앰�\A~�� ��h��e�[�j�;�8a����k�?�5O��������͜����cO@�l�ělIhU�.e�2�5q�Hi�w�� ����iG|�y����oMͰ�9�<5����i��J U��G�;$`����J���i�]��� ij��s������ć����!0 e�0j�G�k�:)0�
�LV��AY?(8�_`�ۥH&Rz��)Rpr��,�Ծ��BR�~(��<�/��, �Z���3�6yw��Ҹ�$r����+csJ��6ަ>�+eJ����y� ��VjOK��n�9n���S:��;t&��_��d삐1��w���놵�N"�kVJV]�e.XwMp�wP�)=��`"���ܫ��[_#J�ԐX	��Tݑ0U����f�S�i̬�4[��1hVqi���*�y8�{���^�FlUGtKLp�u.9)����B�S�O�����#N}��Z��Q�
�p�'o�5K���>��� (/l��
��e3l��F{����1x�tVK���ku�X�C!\�8�>&�!~�<2�)�1�|a�8��������d�lk�}��B�zF��bF7�_��rbe��>�!��|��9���l�em̸�/d�ʈr1��ǎ��d;]�*�[J�m�q_]�pv���46���-���r��Q�b�DF���W�)������#�4R�&�s*l/Җy~�?��=L��t�t���3n����^׍B�5��~�����ΆPG�Am� �kI
�k}i��kŀ8N��Xme�����)�����rQ��X��+@/8�r�>jx p���\D'u,`0��Z����W��b<�,���U��&�ƕ�ȩ)q�3wZzT6���6x-��J�>Q��w���3�<��tl>�<���>ݳE��� �TT����j��c��r�ș[�=_E�*l�������i���R�zl N7�._ӆ���[��T�,�����
t���MqL������%�]t�D�l�(Dc�J�������`1z���L���s�"9��J^�٦c�C
l�7�(���nd2���J}8���HL���TC0A[+z�V���$�[ǫ$�GSa�/�I���?��"}��\T"�.J��Íw�)�>����.���j�`�,&���T�3K�	��yP��)-���Jw=jW)�GS�`Xl42)k���ش���ء���;�ri�6"�~u�� 7���')`Ü��ϒ>��{M���^��6�����(�:��ӷCeP�\������ӤF_#"�xd���� Y$@�]�m��Bȸג{���4�+����R~[���)����w�� �׍5�s�6[�M����j���"ʲ�2���m���/�����Z���_�@ˢ�Pe�ly�V��w�x�&���D�>=�#+���ޥ뽤0��z���<Ad�0�o�CE2W�"�fq٦I��l�t<��K�]�⭇��t��A�'!�����*��/~JCy�à�Fe�-�)��O��n�4��}�E 0o�B��h_��!��a1?s�@X�Q��-k��ui4��^8v��G��0�aY}�F.ܰ�p��\��ꜻ�s��-T3�� s`gF�5��tfE����fl0LC�m�i^|%� |��4��E��g�^�GR�+��O[����F����;���_¿{pᗘ�"�]o�w�B��:;�(���z�d(j�e�a@H��(;�����8 l���ޛL"5�c�fy8��(��.B�D�X�]5���A8��Y
s&�h^^�%I��bC|�v��?�xo��s0bLv���@
BK��{j_�RBV�EW6��t�2Kw=��%h��a����	���pٚ�y��� �Ò���'w~�_�V��T�0�5��wD:�XX����'�\u]��h��lδ`���E���A�'�ؗͅ�gF1!���C���>��c.�:�,���k����r��J6��2
�\���}nP�x�,RwS�T/O-]�ۅ09����s,9o/1�>��9Z��2n��3���8�mȊ�U����JmB_c����T�����Or����,���eT?f*��� ��h�G���2�3��Ƀh��
�8�}��kH���;����B��C:3���\��	!�/2����o���G'f_��S?��Qk���C!��n�bF� ��y(d�Y�X'�q�bg&�];[U�g �}bF�#�A@b��+�);�pp,L2~f�e��H#��%ϛ8�AQ�FC�����A\�xxoYXgX<���[Q�M����st��CfF�ϩ$� ��~uS���̞\���p�G����b�������
ҥ�9����Ab U��V�[�Sr���k�=���	>E����+],�d�N�u��Rg��ϧZX=�D�����v�p4���Js��H��
)�����0�4���΢P�j�x���q�y�	5
B�L	��={U�[e�Iu��ee��8�-$��y�i:޲���Pg���|ˑ���>�!H�$!V.\�@*D�ˑ����t��|ş�r+����I�ya�p�p��RMGτL������5�k�xv#�U��(!��v�z��X�I�Z+�����v���Y�0�ډ�?�w�5��|��.�B�e�~d�×62�9na�0��&c��s��uR��^V։�hq����{����ӏf�n�%9.H��M}��2�֖@39L'�Qِ��(���?`8����h͘x��V׍u�v�c�]���Ae"z(H�K�h^�d�_D{�b3K�
޲+�<�tp?�y���&�����x�]T�俺GI��W�:P�|�bY.*v�p惢��VƱ7]�J�@��I�Tk�!��*�c��ϓ��|rN��������#���T�7�(N2�>���!��2q�c��l/��[) �����P/u��d��M����'<��*�)w�A�k�.�~M)��<�JZS�F��C� 1��A7�/WYp�[�����OnT+I]�(ј��{jf�,C4�f�t=�g*�.�#QCђV���u6���６�=��j_t1G��y�o/r)�M�N��Y	��0[fa�g*T��r'oi�������/��!�W9���:���H���$��V#  ��#���٭[�W���5���Tx]|��e��8���TwYՉ�g��(��� E��f��l�%^�S˂9�3��wj#��lA?"+:h/uo(��Q�mІ:��R�,qm�}�6<Ә��6T��W�| ��B�?��&�ʷ��w�z�]�4'���7���{���7���.Wq��5ϰ.J�� �`z66�������I�h�l�Z��=V��Uf4���o�#t�~����"��<��sE�(		����ڔ�J�o��?��Z���naa[��9�k���;��+m���Aꞛ��6��Y_��~�x��e��b��/P;�9�,��NE��\U@�81�Zj�]�Ҫ-�\���_]���4�d�{4'"��y�>��]R��dMg�#:f�%FcQ�dv�F���ˆ8O+e�o�BM)�:�4��fcz����X6s��ֽL�{*zQ��&�}�(�$ 1rw�"�}���if�k{ڜ�%�%���Nr�/Xs�U>Y����f:'��R�\P�Y���}�
�U���yUb���n�L�ߙ�Ի��wg��	������K��҈ݑ�-��c*��U*zQ��8l��)a�QY�%E͇�5�3Qp���BN᜖���^��]|��	ؙ�u0��=ob�|�1�!����!j��Z���)�݅ep���K~%b.C�	�9���0O5� �j�4=��Sa1����8Ж�a5�D��KBy;�7"c;}�v�*m�՟_�?F��%b�t�� ��F��O�����p�yyl�&��#L"F�:>�&[䐱�O���Y
�KN��p�c���M��*w29�f��;�oL�?͒�5$��f����~�H5���v�tj���Ѱ&U�K����U�%�����	$�j[��C)��^�|���>X��Xv�i��sCY��\j�Vh5%�Q�	����c��$n|%�I��`r�,��B�G�(6�L��b��B�\�q��,Z.�7��c�8jx�CE������y�^�*�̲&`��o�p:��Kl��#(��\幑鳼+���$%�N;�˃XU�2�/YG���ƞ�	J�?3tE����Zu��>d��m0X�c�Y���n��
KwrW������G���Y���"�m��K�UU�O^�C6k
#�� ������8�#�U�Z5g:}���aA=��!/!$ά�b�#�����&��A�P�� ���^$��7�#�S�r��:�h�-���(�����nFB����>�r�B=O�&�t;_��-��Y�o�|���o~:�z��v����ed����N�^�E�:�S��i���V�t{�� 9����#�i<k�
��!�i� ��XgJ؆�V �we���g$̴�z����P�8�2a�>vIa7�
ͽ�k���&1e�� ǘ5=�T��z���^� �@�*���d��٘��H�����O@������m�+4\�O����>�&`M�!��(&������;��ӛ��1�n�'�(��IM*W"�Aҙ�9n[u�]�Y�%���5x.Uc/��df��r.[�&Ho}��	�ퟑ۶�2&�M��
U�X�����5y��P
R���(1�.FT X�%��Z��@5n�j�h��΢ɨf��Y�dR�~��@��d�ߣ��lu�U0�@�	�R�dOX�JP�	��ط��޿p���^�3Һgj�cZ)��W����� p�v$�$���>�Qr�#v���9J�}�yx�:P�<D�x�m&A��c�q;*��Y��?I��e�pg����}U�Hͱ�W̓I�@�:�>i
�ZO~$�B&X����;�H�5'�K�#go�n=�I����6�Ѹf�ڮ����Y��_*�h�"��z�N�s'Y,���!&[���+,f���ٝ{������o�Ȓ��Û�&-8��ǵL��V-�Z�Q�=w�|���y��?&�{�3^����8��T�\���S���C��6}T�g��	�5t�,�� P��Q��H(���V�����e�7�*-]\�g�k#�~� �ŧ�#]�\���$o|q����(�"/�����R'����9�Q���uy�O廵,�GV�����T>rϐ��[���A���(V+n@qq��L���į�8�n7�P5PdFR�>��}0D\k�=q*����r;�u�x����屷)�:N.)ٮ1�K�ݞ��A 7M� d���x����B�g�Ee(�� �/��&��_rf��`{�Ŝ��+�/�و6k�A�[�3�Y{91���| ʼ���p�]p/I���疎�.^��V��7��w�d�>Yd��^��I�����'e�ϥ2ʗڊV��
a�MD�b�$�9Cp){�M��{#{��ؔ�^�=oE�}��Ѭ�Mg�����p�&t��ƴ��E�F��K.�<$��s<F�nJ��&}�݆���a���Q�������#h��䙀�AW�J���ɵ����s�[I;q��7����%���b�����[� X��2
�Ϳi�+�+(72��mdn¯���B�R�|���`#b�L���l|��0��[$	�m��v�t��0�sv���Kn/��X�wE���L�;��D�2��s_�%�ywXܬ�x?�$��I��j��#t{�|^�EP��=���,d9�]�܁^!�:5/�!,߮���T=���Cx���*�V(��
�
 �1c91���,���`	�"{�/8�
"�B��5:@�D��|a�ԣ����h��u#o8Y;Ʌgx��0�.���^���z|� �nȞ��a��/�'��p?X�s:���(��,��Ì�fD9���d8�ݜ��QL��$���OE�ЄMH0h;݉l}��7:c,�0����^��hg��#ΠiA���E�h"�U�p����8,W�3g?iN�9�D��}���*�����؆�Α�!۝�&"�W��§o�
��XV�~�E���rDr���>�\��j��
���x�{ӑ�@a.�n\e�����SDw?V��(�d�_�ٝ���J�G����{Ʌ,T��c�6������]褒�7��@K�R�>L*u���H�ᒾ毱(�퐦�/ͽ�wVvT�ң>�kbP	�쬁��P�/o,Q9r?-JmjpM)U�����:��|�ԑ�����dV1B�K�ם�35�.�ι���8��-/��!�BCm��`\sQ_`H�GƺH��R�؍W�l0����!�`�����πL��q��$�m�TX�!�8��]o)�({^�b����-���믩ZIc7��B�ť�Y�7��ۑ{8"��������7��%���1��,�� �d�9��� .Y�]V:
��}^�i{|6�7fw�Z؇��C:&[1��i1SM�V�P'Ïc8F�=��]�	u^�EC�3.4��nZ{ ����j��_��{�:HO�qx�HG\�7Ԇ�	B�Z�3�����h<
D\Z�Oޯ�_1�.f��T��yu�[�8���hO��r$��E8�w�5,M�Ps?\r-��x;�YA���Q���S�b_���n��%�E�\�/)�grR����\��+i�7�F.m���ݼ�&ʩ�v�.k�"�}�����.��$x}�Z��k����ۉ����KfW*2㖙�"ݏV�`�7ƛ����ʣ�����R�q�̌��z�9.e݇܆���.�8�x���|�b�f�,P,��rɲ5P�	'��:�'�߼ZB�x�o��/���͗�� ���:}x����)WbW�^��c\���{�8dK�8A�XK�)3�":=R��L�wW�g0�	��'�-��W{��|I;������>9ۏj��0j`����C�ĩVH��w��d�E����m$�F��,Q���`a��+0���@p��t�۩���z-��%�V�Z�̸�$�M#$�S��z�Hԅ*��ܽ �ܖ�+%�,��le;��rj�g�{�X��Ɏ���r�k!�|��tm�`s�	��<p��ڨh0����ur����/�6��O��2�j�|ݡ\�p�fqw<c>3BL�2fԌ(;��dF�zֽ8p��=j7�����<��)�,�K��W���*�C�H�i�?��˭������p.�UL#
lQUo޷v�g����2%)�q2���J0e�g���?S�sS����щz@��eZ��k�tA����)F�,\�������+ԡ�d`a�r��l
/S)���K���@n���r����W3�(�6��3�j�\�����
q-~Cd��]aN�����܁WI=RO�aN�ت���Yf��HL� ���Evy�S"$����헧^.�����Itq�i�Q��T����̻�h�@����z%3��A�n]�8jU��f�<�2�����Ų�����x7�����mB��桗�_~3U4.󅠱	GfDv������,�X��?~��`q���bx�Q����M"ź=�[_2\�P���]���5w�5��E��Ɏ����;F�-�ɿ)4t����(��ڶ�U�I�SC8�����#�&�����<�-'i����J�����
�wa~nO�She�g�@�:v]gz��� ���m��|i���Ak�*U,N31ޫX���纶r��a�-�')|)0m��92���"��`'�Y�,]P�m�ہ��7t�YX�R��d�f�Þ��[�&܃�8f\�X`U��u=�h/�ښh�F����v��S��o�fD���b�O�j�3,/�,`�#}׃�k��U�щl>J ��E/�\�����ʩ*��S��Ě��z;�lJ%_�w���ސZ�13�T�|_4��(�l8��Ќ�w���PrD��~4�i&�蜡�o�u��*B2� ��Q&��K\��`B�V~<ç�r��ЛB}Z��mf���e��B4�{�"���LN�c�+_�s��k5.�;�ώH����Qd��9����>�?p��^Z��i�j��!'K�q���o�<�!�$wm�!
�,�x�s�i�N�f�Ն�ݢ�� ���e[�W[sV`�<a��\�SĸX���mLrP���#t_�z�n�#�YIh Z��Ƈ��& �aI.Aُ7�%s���������@T���b�5~c�)ʝ���YϓX�K�}���!�k�?��ɡx����1��쓷�|�@�w���b�G�YW �au�΋�$�W�Q�i&~4�٩T��j�{�pq��@�<��bJa+O刲�:���V�Wفn��cHB��ȼ�������.zk��(rx�SZX�wE�����50����14ڣ�}	g6��z�o�y]H
_Y+��� ?e������:��ai~~5Uyrh<Ѧ�� -��lO]D�2�lCd5/;��)�m���$�G�pu�b���=�	�	:���I�LK��yЌoD�|=D�²x��ͫ�s�R?J�+F&r`���S��$>���e���0|Ѷ뙃���Y;5��I�Ȃ�w�5W93���#4&ᐾ9���.����h����mO;�g�3K8�U�y%������b�!h��#�m���<bv��Wk*�C��l�婸f_���:G|c���@�{�aL_�wBV9oMڡ�P�C�og�'�mj9 ��jEI!&cz�I��n��|���y�O?��⋴��Ne�ca����\���c�Y��7��)�d����~�R�l��E���t�=�5!�1I�T6���dGA�_鏌蕘[I[�d^L�5[Jf��۱���<o����R@G�BK�|�<P�X�3���k��	��ȃ�^�
y��O�>�`�ږ�rh��p�'������� ���L���J:��GWJm�;%q���_�F=;UBa��c��H�jPew��{�����#e�Z=9wA;4&��;6�	�N�8�ޡr5�S{ �v��ó�TN��1��Fb����f�'R�e��Pw7�֠�w���׼w	b!�cޞeu�7V��`\I�ɢ8��D�<֦E�7�l[�o��v�~Dn�l8�5d-Qw�O�a�8���Ŧ��x����_>�Z���H�!�ufQ�Ҫ�,P;j"�V���������!ӫf|�6����	��7f�WxM\7m���Q�љ��/k2�>,� ���О!�&ߤ*1<�������)B�����%Y����9#���]u��w����ڈd=�^�P_zT'�5�(������-
�����	2�p�Ǧ|��'�n�9d�ل�Aw  ֠�D5*�!�^c;I6�bo� C_wj��Ү�m�������P���Ź; �k#]����I߀:Z�v"��ԛv��R=@L�O%�b�(ҷˈ�8�Z��@{�-p��J�0ٕ��Ȥ�57]bl�2�Z��eW#�� �Sj��u�A���z�Lϲ��(-���4��퍺�̖�ҽ��8xN%S�������V2C��� �1��%�门�$�L?U�£����q菕��Jym�'�6�=�Y1ٔ��N�����	��B	���{1�*'�^$�{|��ߔ�w�S3���<]�-Y��|�/���s_���o��)�<����1�j����fN3�i7��:s�L�M��@���Cś�<�̙Lh�M�FeU��~��v�\��8md�� �2�B�)WI7$�sR��8J�-a����U|�	N`q#@$j�)C�O1��+�H�wz�!����ǲD�R\і/��c?U�,����}�4����[ʢP����Yw'��ۻ���Is"��|��h��r:_9f�Rg3���'�W�a��Y�vn&"|������հ�R�I�2�bڑpC1��������5�^>(0M.���;��>zy�I��<�/w�<rk���t����̿󟪱�#��+� �la�r�i�S�COY���lFA�`и�.�p�D5���>�b�Sŋmf\7W�b>��e}��Y�W�������W���lJ��9.5
��/L�A��!�.�qu}�|���|��p�����so'��	�Z��N\��ΏV�"y]�lZ[�z0ՙ��4�O4��;8IfU����dCycv�>�����{7������!�N�������H2!hV���!���|��w
���-V��J��H�[a|ܦx#i)����s�>�n7��j��.�}K�dG!@?��Z�~� 		��)%^� \� Ed�,�{	{6y:���޷keц����M 8b�Èc���R[�!�=S8D"7��Y��$�#6�*呈t�G ���t�
�O{	�~��2�T���Hy����q���+ŏ�\�7�~��:��u�������^چ�H��r�GIv �-��֨�(�'�!%l�<�ʄ�=Ch��yc��O,��r�0Ի�撳Ju�t��<7��HK�T!I)��~�B���	�Ђ`E����h��0�T�U2?.��о�R>��?s������F�KTF��s����^���V5�[^- ��u��9L�ZV�2� �H[о��ܲa�<�hӝ�BuLdͩ�H���}P_�`�L���[O>X��$$��.�Sv:}��b5��:4����1�J�ܾ�����Mg����u�i���u4��n���	�cJ )+X�-�A���(0�d�17M����xi%s�-c&^ޥ���W��	��6�U�T{�s(C~��+	�h�X/6׿�y�7����-Uʮ�|��,7!XYH[W<>S��DhsT������ے[|>�D��a��M��//��ň�&Y��8	�
p�~��kk�GԾsP�!�"[p��x1ՙE�!̀��1��2��$�S�AX�NSǯ9��k��u1��C����?1���5*�����¿]Pi�g�)�䛧ŷ�����%��z4_i�+�ߧ;f@�[���7�����$��A3����"$��\͏_G2�"�E	�;�@l8�@4���@�_*�-�>�PI��x���Yi����ڴ���k�4�$�d�����~�&��)DH�����'.!!5�C��f�;͹:�ߥ����|\o�95�.#���隗ò̂�d�� LW[k��ev��P�
�\h��#�<N�z�,w �>u�kǘ�j�b� ȸ(<|
��>���F|B��)���*"�����I���@�|obh�Ñ�<�<`���Ʃ��p��O�RZ�?�A�.��� ��vY�S���M5��6�rF���'za���w�y�`Z�iJ�Cei�4@r1�V�j�p�a��A�v�Ǯk�^<$Q����T+�p\c������;����_���l���<�(�KDT�-�+\O�С�[�|o>����8sE�i2��b[�j�S٢� h�����Ό�mj�p�I��=;u��u��e�W��z�����rݫo�mzTN �}��)�d�R�K�|��ŏ��l)eJ��c��,�� �Z�yo3�+�P���*K�S�S~����h���v۠}.��2E�����������m(/m��ͳnԥ�G�s@����̽=��Q�f�ǣ�s�YkXzү�ƥ����TćQ]>ܼ�lF �/�{T��v��5#����L�F�y������a�}��;��e�nȰ[D�6y�͹�_'w��!�!�y%�)xM6�`}�M��mb
�ã$e���ʧ�+��F��|4�&��k5�6Ǡ��o��>,$S�v�94�>ԛ�,�����s��	�`&��T����#�!�˲3Y0*��8�'������V-w5�
tˁ�����DȠ��S�.!���CS��J;/�x�0u��&�yB�G��`^�X򁝌}�� �s�:�=�y*FFGvNt�H��UgZ2���z��V<G&��v�I!�*�7�u�|{�^B	EЂ2��n8_�)�{-x*���E�M��_�bcƹ��6JH�=9X~����<{dJ��0����Ji�Cݭ��_�������j�W��u݅��x��`��箴�N.��%�t�� 䒴L~�Q����r*�MA6�Dŏ�����o�p����e�7A��ݺ��S��V
��9͖z�mAHZ����4<*m�h]��ȟ����N6L����|a�\V	�������|[���F1�ck�����(#���m��$;N��޺&�,���{zu�u��A�n��s���?�:�>s>S����r�,��
�)C�R��T4���M�6
��>���#�6/��e�'-����$���.]���[}ˍ?F@6�3�4��T�b(�{��Q A I,:Bd;��t��;p4n�a�O��=ړ�P�p/�$�-�[���jS=�1��Û�d3�N'�C!J��w�f�7b�N�"B���¼3P��~�����0 o�ÿ�nTX)�N�Z���/G�K��VX���>��e4�R8�y໖�}�ɾ}N�m����,�:�=�qA�X���aHY�%�)�=���g�'_%���j���5�\8�]sbbI�JOM$�;�v1B����3>Y���$�G��x���%�˫<2;�&�v�%�/�ۗ\�b��hlŇd`k��<N��0'
��;�����\h��fr(7��C�I�~O��A�`�z�א�9`)P�&��Z.���ڕ������	@��sݹ����餾���
pu|��'qgƬHgI-O�%%��C"Ј����#dKu|��f��_^؉~��Dj�?pЗ��3�Ѿ�w/�w�Ԥqd���s�����˷�ͽ��Ʈ�3(��G.]OO����r�R�@��
.��}� �C	\��bQ����k}����&�����@���QH�z�o!gI���;�uo�);�2\@��D��W�A��ME^6���W�Ci׭G�����/��j�8
 	��}>R�(W�8�f���E���'�[$J�?�,�Q��<�э0\ʺ*���K:8}�_"�����vUe�tIwS��vY�I)�	t��ݷ��s(�''��s�n�t^)R�i̤�;J���#�F�̞�;�����^��vo�2 ���Fƍ�=\����o�X�����j��&�n(,��ڮ�z� �����Z�).d�.5�fl@	��O�n:���r�y���bDq��Vi��=6S/�@���a�>2]zd
�4�F����Ǒ�<�h��ϩ�fc೦�W�7���q���c��t���?e��$�R��nJ�~���_g�&��Tp��kԒ~E�!=�H4Et�,x��
;��"6��������(��{7�R���ˑ�0��몐Y�8�8�Ʌ����6c��:RG"�֞:�WM�c�p�Vh�Um�7���Nڷ��F�"�T*�	̃��K�h$;m���b�YH�}Y����m�a�JM_G�����!P��]?cr��U{�9����.고�r#�ԩ:w{N�P=���Λn1��+ŕ��"!�8,��N� �����9��9O��oM�'�n�X_��kqjBɺ,I�QaZ�W�WHځG����BG��[ic/�u�m��d�4���ԏ������S���������ҵX[B��t�2�3J�J�}!F=
�r�)M��㠌*��t�sGB[x�,�P�/�聓c��R��%�'Cƻ��w�<<y��n6
֤������r�1A'�pI�
tIR9`�<��E&�`.w���Vח���^}xGm��ƛ���3��~�{��0Ԟ��ҁ�:�&�9'*�bq⍗�Y�eRїL%�2�	���*�<�9�(&bRLq8��?�H�^r�R� n���B�C��U���t��G"]9hr���o�t �v`QL���9g��\m5�R���b-VIJQF"�=G�vV�y�y���Y"O�Ԁ��X�����A�^=����x�1��#_p	T������4d�e؊����-G�TT �\bU�ڟ��<�M�NHh�}G�f�yI�W�</s���PA �
�H ��<�G�����˄�r�՘�BV�>�@��0�m%���J�O��c{���
޴��S�oYey�\�E���Zު�2�xju��K��h.�)��)��t�?��2�`�\U�錒�
����"DiѫF�ڏT����	�����SZ���G���v�70�_LF�Rjw�2xR���O��M|ڡ �Ws�S�Vr'tL��\���Q������sS�c���TYuj�g��d،�\����Qd}�4�z�� $��R�_�h���)��*@/���x�R����s�e��";=���i�w8w��뇌��6�UUB�Х�H�U��Lx�X�r@�|��fd����0<^w0�v8?vIOK�*f��k�a��Hz��R�N��q\�ۼJ�� q�ڃ������R��d��4so)��'���q��>揂�P�s�c�?���t� ax��hS�KP��<��u����!��}"��vR�Y1���Dg�]D��[�����'A�Li�<�C(gfv�O	��O�������,��3���i�wܷ�������LC|�ŤFti�Kdfo��� �T5�}�6X���#��=vP�m��+� Ѣ	W��ٚ�}̸]r��f�N������/���Y*�V����iM���VW^w7�7NB��$���dr/��p��4��M!��|�8�-��3���Q(M�׉��R��2OGڗ�P�����m����@ڰ��/��HF2��b��(���O) �*���ǣ���sSf?�$O��e�8�|	`D	ğ������5/��v*v0��\@��g�}i�]���w�����-^�Q��º�����4��0a����q��?�N�p$��G)�i��u���`Qdke�?��e����Gsĝ\�m�A]�愁B�
n7�p�k���;����V��cN�4���I3�"�����a���+2���<��M}��yS��t�gP�7��#2:�D�X��Eȳ��w��*
���e:��q��a���IB�S Z؅����a�����'�O`��\Y���������*�.���)�'�L>r��y\��t'��t9yvB�k��c�2oq�-_�v�����9H��D�f1&�����u�g<B�ꢈ��c��5�\�T��BlR5�ּz�$	�qH�+���P�ΗD���d��Uf|�z�������XLf�Ժ�ha
4uXA���
lMVa3��Ź�*3$a0����_�*y��R��s�|�`=���$
c�>��	,P�&�{�z �k�\[͕����1�Xh�b[C~�L���g]���cF���H���L�?��4���ؚʳ���➉M�v��Z��t/��/s�����".l��x��W���dRǔ)�����*��u���T)�ϡt�~H�R�13s�,4������MA#}���^�	�~��(��bN;�"�����ă�0	
�Q�m�UΡ2ソB󠙓��I}� ��`�tB���՘��~$t*��\�r�Z>�z�* d�+>�E��O��a�*��d���B�8	|i��%*)y|����-�+f5�ʦH��M�<#U�n�/��6�6��)9T���/�.w��E�4�E�	5zH��ɩv� �~4��� �IC������zg�ي�X����KE����M��dE)��4"~iō�91�Bi�OJ ��O)�װV?:���*�u�Y�;k����
\>���t?/8{PQ#ʺ�D�зV��ҦU���4;�m�f��c���z��]Y)�8(ƿX�dD/uYt`3��S�6�dFT���|0��XzFM�G�@V��9)���{Y��ZA��@NP�]�DV�b�[u�[�g)���14���jN��[�"}���5ߪ�`7`v�Ɯ�N���cZ݃D�b+�뛫b���vy=d��Hq�T�w�������\�t���Z�f���:j� ����'���i��:�4E�n�<�
"G����psAC �X�*ʓl�F��RfXC)"hJ�Q�������.R&H/�]�tTX��c>G���&��t�Bl�� w���+K�gP�2�
�y��L���ZO�~�5��[5tɁ����p_>�$�Ҩ9Fv-���5q�J	ua�W�+"�.k�=?� �>����Y�dz�Y&7n�*�����TҜ�`�Ϛ��,��퇅I�٪��+L�$���^�*�#z�2��� #�x���7��!@�v���7�Mo����)��k�D�)�`�lP�a��z�t�a��Q����8��Ķ�pn�g~7|]�9mZO��`^����iJ�t<^��$�jJ�?F>d;����e��G��!�d|P�_���a[�^4��z�ՠP�0Sf���t�'��1��в`��Hn�L��Z���+X!�$�{�9�R� N�7��y��oK�4�|Ե�O>U��e}t���4�AQ�N�p��j�u�a^T��pM��T�x��������
�/�ꏆHs}��}�U�td*3��'Mh�l{��A�a���w�,C)B{@��9�L��W}��%��gD�6�V�/�oG3������� |fO��=�,<)��0�Cޯ�5��8�_/	�YD�$�W>�s�p/�Pnu��@z�[�p���	�3�ܫ"ۨ]�c3�xYC���_P N�$>�m��\���K-R��2�mT�~���?��n
8N9�L��I^eQ�&��y��$�M(����.M�5^�iy�s�������*�O��T貘O���A�u�
W-��6�uc����3��/)g�f%ľ��Lp� ΃�s.Wk}C����z�(m��[Q|q
���l�Ixk��yP��+�r�7��Z��+<��, �P�	p�@��h���)zYmY�`M���jBC�Xh�9����+Y*��7����"-���1n?~�J�nmT�����ͦ�6��wE��r�Q$-yzˏw�꬜�t�c�G�5w��ZJ�g*��`EP�����W�x���,#��c�b@��[��ߞ�x%����~&� ��#񡺢��8q~�<j�v.��[�ī�c�OK�Y��WϹ�O��+ �;��˯u��-e/
=�"�'�[-1�p���ښ�����R(�I���t�s=FwC�_d�0r)c8b�B��y��S?»�6&,���<2V.H=k"�+�5� D/�= �"�����z�C���zӇO��U)�������v&x�OW1Ѐ`ط�n��D��旚����"�����եO| ���7�(g|w��s����p�Ԭ����[�`��*����{H�k�J&泿���j���'`k&D�ŒQ��u��#�4�����*��]����mm{�T������ygU����Y�W������N�ko�_!�=�P-�Y�L��d?z� �'^���p����!D�t��K��'<�K�\`%�.�b�=�sݘ8����p�o�(!�O�l$wE-�6�i�D�kE�VX�
r.Vt�\���Yٕ�+c�٪,�s^���;:�9��t�H�rf6�� �õmr?�ӹy­R���?-��������L:�q�ĉ?������|*;�Z�ɗ��a9����F��������G��L	xh����y�'���=�'�0�e0hO���<�:�y�oQX�%J{~���Xj=f��8q@W�AS�ɭ,��T�Z�x��d��ߝ�YV��F�ʖ�"� K��.�<e�Ӧ� �x�J�I��2�e{?�gZ*��9Z�-P�F_�]xMW�v���{�������^n �,��كM6�b�֖�46v�O�Z�,^Ν�9��F�4��Hp��z��-'6v�`WdK�7"��)�u���H�q��w��QIx��-�o������Ҩ���E�#	���%����� <�v�2��x����������pהk�u����� �|Y�)�(�|{���=�9���eJ����4��+�!���|��/�����Mߠ��G4}k�S�4>���[Z˯\K�r�(pl�`�u۔+�9G�-�0>Vr瘵����M�x���˰�O"Ή�1=uK�W�`���6ޔ�{w0�3������p��WhV@����˼Q�=����T��A ��(�#�C��Hu�8p��f{Bpp�]*2�x1z����`+ޑ�E"���IbGa�f_�Vs������*��ϱ���ļ��f2;��^������Fl���Đ�����NbBibފ:^I�P/F(c��S������e�VO���`rr���KV]q��'�~�e,˖ȏ����;}��p�Wʁ�E��%!wD]����j�E_���N�R ��J��HYTc0e{*��ﺖ1����(�8��,�\�����/p�a�?M���*=ϊ9K�T�r�	ݗ/zu�OL���,��/'d2+�f�`p4���_C�|B��3��1�r�Ge�������'�@aK���?�cy�<���q>��h;��48�:F���YD%��2���+���6�p���<H��������9������|p"ك:ۅ�z�g�#Y��1���k�]+�f�?�ܧ�ɕ{�-�w�^�wO^�kֽ>�jɣ��E�����b�8w"=����!�����?� �7�MO[˓w>�*��֦�d�Kk0��tDSe�%@`���.=�r��"��/u}6a����J�����&�tx�ϱiȕzV�)ctҌF�^�n=��ȃ����;��2�/"��2��C` ͪ�X���j�r!�7C��LԔu_�M�Ț}5Z��ߣXlc�r��Ł�����Wq  �U��) �X��?Gѭ9���y3N��E6��b��G����h�������fW��5�Us�cÖ �,0���]@�mG���iZ��L7u��p����?� 8�K�۲~Q ��ciX��^Cc�|���C���^�Ngcb��<�YOQ(�c�)߂�������贂_�����ʦ"}��ѱ��8>fG�J��;V�P�K�D�]��A;�	�yLQP���>D7q!���'Տ�hA��_ ߳��D�@��{q�:w���{��_����vw��pM�8zE\k�_�N���_�Z!�Z�mV���zŽI\lW�:L�~�q�(ǫ'�jG��-�����v��G���N�0c���}*7�}�r��]����
�oA�(T�2��[��rZt���,��K��j�����ԻE�"����O�\���[E�3'�����+��^Y�)Me���`´
�'9M�Z:�b���93���ʠ�U#K��&��G��;iSw��sǺ�E�>���^�*,%)�|Y�Z�eU:h=�{�;E� �$�<I��\����jD���Z�^���[��#�v���f8U/h,���.�O]Aߚ�^1��W�MjZ�yЉ�x|���-x���mp�s���e*�E^� ��(V��h�e7!7F����-5��ܩ2�L��~��'�#���r�dDC��cA�[hK��C��������ꢳS?���OZǴ��%(��c��o)_(ɧ3(�h��۾gU����W� `�\rV���0����*�	���e�v[�r�AX'�F[���p��2�}7�V��(F��I	޾�}���i��a�I%��t@�����qa�W���~��~�������R� ���g5��CKz�Тu���z�� h�`&^iԎ���¤��xTfF�W��z�s�V�5�A� ���:Ҳ9�A�tkƔ;����(h��y��UR�W�iy�/����}�u|i��\���5 �n^���X6������ߝ�?�wЩ�u�^ꎨ��ܙ3 �S�]����{�K�o4R��[��K��Z�[�B�RV�t'�b�^�RN"CŁ4+?D�y�_]�֗�M8�:I�Z�$�R�� ����C���x��K}���s����r4eB]����������,w5�;J�v���;6�dm;9J�BA?6�^
��Oy��\!�i��őh�F/W�R�f���c�-@���lTE�jph�h�\�P>�Xe.6�J���u�7���y)*K���(������Uع�Ð��{�������%_���7(�� dE�4��ixdC\��N�Z�a1!�@����`}:�+��c��L�</��ؼS�����ķ&w!�Մx$-�0P(�Ӈ&�젥i�\�y��p�Ͻ���B��D6��d��[�x�+]�����+�e#I���\����