��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR���[{�T���CK��TC,���:�
&��d!��]9�'D`�"9 S%�aQ�`!�6������V�W�l�a锦E(�\gC�slu�4U5=1�N�m��l�9ў��P���B�@+yg��=�}|֦���ָJ������4%o�F�5@�P�3"W%�/��X��A�JN��{�q�4�ug��H"ߴimN"�t}��-�4~�#3]=��"-~�3��{d�4��#s�0��t�1Br���%-MG�pL��aɳ���Y,)6��%���g���O��.�z(��f%�w_t�/e����O(��>�ig��/Wl��x	�(�"}�y����\흫���j�ut���]���t9S�$aX�&�:�W�@G|`ID��ˉl�����i��&]��D70H^všR-U�����Q0?Kd���]����ә����d-cre�`:,ي��d ;dn-a�9"���W�7\��z��^��/�����Y6�F�@� 4�raB�4	r�K�=���w"��T�<�a�o�Q��i�B�a�Ύi��v�|ȯ�H�K�ZRj�&]ӎߵ.�}N�x'X���6�.95��<�v�IĎ��2h��T�7�K���Q/M�)뢵�A�[��+*2k�x�����"$�,�P��m�2y�`����n�~���E>]䋜o���?ڪ!̙	�tY���.^.�@v������$7J��+��R������5^�,���1�
;�R ��3uS��K��v̃cY�*��(������Ղ���9h�=�7��G��賓�7J1�i�.�k�ˈ��8��)!�r�S[�ނ"ټ�bE�!�Wx���;�n�����	4:�E�^i�..�J}�֚�l��~mY��~X�t^�'`{ӊy�{ ��S�/k.�"h�����lB�-_.~���9Gڑ�?���%A$F?�:s�f�ߴr�W���h�T���n������9?��v�X6#�GeǮ�P��|.��w��0:�h��c���a����b�7�B;m�pi`�~���1Z�o���xǵ�f�G�f>E��i�8%\�v�� �I߷́mS���S0�n���pg��^���*�sD|�#�L��j1��5g��?w㹜,i��^?��ǚe��ؾlA������p9��&\�8�2��h�܁1�W��y�s[�J�!O6�v�<�>�N�㩦��7��l�i���-e�g�]�~�LE.\��bL��Jb+��V/�����&*qxAjm���%���k��"����I=�X0L7Z~��$"ߪ�O��	ϰ7#��3���0)~�L��F�L'�U�Ϲ\�����b0K0꼏c���Ԩ8��7�j]�Lq�����|i2XI�AKCg[�À�z�;�FXySEߣ�W��I���{���b���>�����C���ԕʇ�a�f20���W�!��Q�����y�RVLO������qO�Iu^hEb#��*��Ӫ��5^�;�dsr���Ȝn�&&��Q��FU>�獍�v�2�Z��v���Hߎ��Cs% �a�b�˽#k�ي���:��͌������J8�XK�'�;��[7od���h�����{]�M���)%��@�ߒ��Z��@�F'��%����j^mw/#H�}M��pZ6Kj�Ƽ[��_���P�����]��{J�CU��vk�THV!`9Jml�#Ʀ}� �U�����Xě�u�o|�9?�;^�;�t��F	 !��?���Wt�a��� ��R������#yj�����9J.1
鞈�����;$���?3�'�0����X��������nfC�ۿ���қ��q6�O�K��A5%6�Zq'sͼ*&)L�tCP��<�A��G0�1��F�h��V"��8�c*��_��ד�K�!2�7��K�^0���پ3UB<�U���XG���΁{�wr�nzL�Ac���&�Wmk�,��23�&�r�M)��/Q�2�	fC I�@��>�s���v��22#��k�Oϴ�
��<�0,v����_�#�����?~�����n 4��p�4�qX>p�$�A�/�-�1����yK:έ�=��9ձ/��8jF�W�T �<�'�[���i�aZ'�>��8��G����F�@��k\b�eo�Jr)������$AP�Cן�r����@������+�AY��s�t��6$�4Vdː����u��ɽ�2Oo:�by~���s���)i�I���U��i>�#�׸�6�6t-�����=K�O�Q��hK�f`��[�?�X���-��&����wu��_���j[ͪ�&j�R�J�)K������0`��0��ҵ�Yf��jZkit��Mn���X�F+�$
L|<��dFmBQ����Z��<f��p}t�i�����N�I(xv�|G��1c�S���^���$�,Ejd�y3�m`��w�����6����tB�\�Kwt��w@�O�O?oP�,hҔ�4"P�~K<���#�2��yV���_/��7�6�a;�z�s�dϋ(Z~.� �}yMRR���!�E��{.�U!�tL`��B����0�z��<�m�A��6�,^��E��'��իrߍ�V��a�E����3����/��$��Y�K��:uЎ:�!VI:[@#�0�XX�ː�c���z�^<��l�z��T���Zd��.��T�&?Vj�=v�}�%��Zu	G�>�/*9EN�Q�{�/����`�kt487N��t=3�'w}B�tDa��zr�����WS����g�H������ǎZ�	��,Kq#�~�_� ���8�?��g�a:<��9ȋ���Ns����\+~����f�d(+�%P�*nn�<��2[��˔t$�-�O3.�lx���d/�'xiX�����h���f3{*[��v��O��	���%N�f�L��8;��	E�Κ��b����
�k���ǧ�w2��O+���*0Dzj����A[(�������G�m�����K\G��p��m��g[�����`9d���'ڵ��b�����d���̡I=:;[&�"�V��N���Jk�l;RYN|-�CIPa��!xGDs���54�8kz�VG��t~>�:=s|J�?��g��>��wB�9܇��(��>��@JR�%~oT�=I����l��$gĊ�T_DC����K����yM�zR�H>d���㷤�蔣%�PQ4�ZN�\imkQ��)S�ɕ�?];�����BUjd=#ʰe	�c�$�`�~����t.�s��J�p���頫>�4��7~�N�h����������������_=��H���J�?�y��?���Q�C�w�V�o�*����qh%�����̧��& w��Z�C�(�7bg���t�_ӭo\'���s��h�fl�L'�h8����Z9�H����L���݂C��s�$&��sY�<������������٠ɛ#�ZЀ�f��|��M7E��⟦u;۝_d�8�?�����{�0�O�^m��NE��\&c��o^���ߺxz�u?�cR��{:���v���Np���K���W��# �����t�}(�&��Q�k�k���^
о���'j! ��qp�\/~��R�����67��~[�CZ�"	s�2�x�I�(���k���yj{��(>���*F�B�᲎��C���H꒡������5��p"�4��B��g|��e�P��9@��������ˣ��t�7��C۲3�sw̓�e�-j�q�m=��?mM?�Z��I�9�s��%F�}��iK�W����ʇ��x$|QO����cI/�ᬱ۽�5NUf!O�YX�vop,�Y�8�B�Sލ���'���}�j�j��=�t��6�����.�RӣM|���ύ�Gxۡg\0r�Cp�s _�N��:o�G%a�mz#�?�+�L�ٜ�^p.��p���(�x����g�]��l?^��?����49��o�F��_Y�C�lс/h�GwZ�顉�ma�q	�!��3���ޝ�"ʥ������{	��{v�t�R��*�2@[���� �������T�0@B㱟_UA6������p2�Y��mKq�������1����2��0Ek/-�=����{������0ԧ�8u��@#�됢�?���"�b��n�9�n���J�&�G �fş�eM�O��O�Bi3�P������x�s)��Ѕ�6��-�}��~��8��� ̄#�[ ���M"v7��dͫI5�^�H�,g7�T�����߻�F�2���3Y`!_�������`�y�����f��|�u���ņ�ή"��_T�~���_.�NֵF�bi{��{�:x�c_�6r�ޭrTB�����r��H�.O[�NӉ����'����p>���C��D��I�������1��C^tɽE�mm�DQ�8�Q��6�0P)?%?(��l��[�E��Le\��6���[�H��ِW$���� w��)�����B5��&�y�$0�?0�ů�jkh� j��Ă%�w{~��^u5r#u�"���R5��{�5
���I!�o���h��~[U��+�tX
�tyQ!��h.��֧�S~:��7)�<��P�[D�ms|�F��=/���9�^�~o%�����C֑�-��~������S�EU��P�οѢ�W�����:$X>��~ Ci�Ň�K����ImA�N>RY�Ą�SF����,.�9���*�C~Q�14�P�V8��J�ٟ�56d{��U[����OGx� ���&�o�e��b*qp[b����U����d��"r��93/8%k�mMP�>y]�'�?��\���v�˙��NV5ub��-��5V�,h?�&�+F���"0�~A����[$ͨ'����)�5&DP�12�xQFU�7Wb�Y�	?1�(���:��u��u{�Y�#�Rjҝ��j���$.-3�NȨuj�h���D[!4��yJ�D8�u�'��z�0�ZZ�AL`�
��	�M@H����s��8/v�W������mo/U!'G���T��N�b�[�ω������;�G/UX�\���h1Uʉ<�ᝄ�H��b�A�!gQ�f�C�Ď�X�[ ��K �[Θ����ЛY���t�/��͝��	5��.������.A1b��o7>,�O4�{�:������0�#�d����˝aQ��}�]��A��2[y��j:�r-����'���?���j��|�]�ϧ��i�u����P�9�96� ��_u����*B�D9�� �����i�R�&'$����z�3�R:�p��N��@�ۦ����1�,y���ϳ[��{�A��P�x��J���[ST�9�zّiK�m�|,tU�L>��P�rO��nΦD��tb����7{��A�=����e�i �L��m?\�W� ��'����m�;��bP���	y"�DE��_@�z�ԛ�Ԍ��g�1�T�#�zv���\���;w3o���z����p�v��TΫ�@=�ˋ\�W�=:S6�;6���bR��SӪ9q��E������=D/-�kޛQf�pGg����(�OZ��E�f�1�1�s@&�x��[����IX̋>Q����;�k���=��x���?�FK�o��
�@'�o?�����H!FCl���B G��0=狆<6��0&��	�?�zE���P���-���u9�Q���w9P��5�"W]i�/���K�-�ʵv߶G�8�?bIGM�eo���f�Ƣ�뗼	�I�����>"]tF,k��џ.�-J����K��Y$u�����Xg�Tr��qf��˴z���X��ҧ(�=$���R)��a�H+��5G�C��ȍ_�(z��G�N����V?Vu!�xV������?���
`���X��K��nyg�"�-j�4�_�d�h�Z��h���'̆*��3�s5ȵ��+���]������=A�t�@��ܧ�|0sA�;Nw0<�,=�`�\n�sh t��N�=h����aH�J\I��l�;r��8y�H5)�e�s��)�ŔÆ�^��e覸�~���h�6���<��--�<vuȪ��������a��f������W\��j��\���D��,n'k���2n6�T���w�#oQ'�3�.u?L���k0�e��3M�<]�֜�P��9��f�����Ͻ+�r��>s��O �Cd��h$\ (��|�,}����Y����k��s(��oŮ��-�T��V�.UTE�@/����Ο�&-6��r�e�z�C���&�O�e�\'��$$���������:�� �g�[:h.{���w}�Zp���9D��@g��DQ�~�l��<� [��o K +��5ׄ6�iP��� �DB��� ��##��m.1��>6E�'RTڍz���͸�Bze_���dJ��OS��ɉ���Uj~9s�j�&��U[�xGB\���k�vE��� Խɦ����mݮ�X�_�z��7��I�h��z1kw,�u  ݜ@�d4rf�����̵�O��"ֱ�k�t��.�������ᘩ���2���ш%�ڊ&7Ŵ�B�x��SX���XJ��W�n� �/��R���ѕرW�� �կ���V�K���A��$�D��b��T��Z���`E����}�� ]Ye�;�D	�:��3��n�<��ƹ����>�:��?S�.�>٢�<�����H$�Ogd��x�Xc�T���h��JM��2!Y��z��0 Kベ��î�o���D����ԍ:��!���fk�=������FkB��_~sh�h/��c����rc��˥`�&x�!g9�������c�n �g�v� ���*�N~���5��9��Q�� *jP!�YAi�&�
��YUAX�_��C����Q�J����À�קJ���<�SR���.�P�7}�4k��A.__�s��}����w_��f:��KM,�2!2*����߿x0�u��N�e7}�g�n9�uZf�Z��mtU-w�5���9Jb�/wJ�<2��̥���o���!0��!��T��0�mI?.�ץ��F��p����~7��܀�����/Sg5�#T��l��ض�蓄0�K_�h貝�ҩȽ��,��|�ȯ�H��A��ڻE��Qib�������6���T���_���dy��%z���LE�*�
�@�1i>fkGj538��YE\��R�x�d�$|5��s�0����3Bs:<Q#L7�!��}��'������`��5��hz\�z��^)l��)A�O��U��͚�e���6x��$�l�,A���B�~2��CKm�p�dx溠*��F�Lѱ7�	A!rd�M��Q~��m�6^�_0&0
i6�qo�E�m�ҵ{.�a��.}շ���q��^�/�y�P��T|�}���½�����K�KtT��3�,�7�	|HӜ��s��e�.�=(�ǛN)B	�V���XPlN.�Е?B�-���'n���{��>|�n~?��X/��#*L2k���t���J� ���Ӕ�0/r0d�+}�r��yHO"禺�
H���Z*y���	z ����_�OE�{�/��ᅜ��]���&�"li��pՐd_�"��$(��e��*�ȗUxݤ�ھ�*�h�HY"���,��a�]7�<�M��u3�]H*k}?-O���'��'(^R�^��%�uJ��Q�A�~6^���G�2��8�h��ְ9/٦z̽�[S!�>�M�]!��r���M�~sZ7:<6Z6W/izI��n��]D���ܗ��ê���L���/�����o�/��@ ��+T���}�r zǱΔdI�=��3Z��:���û+[�N<���_YvPd��A�>�e�XO���BGT�slֶ#�'�� ;���-.d_��N��ǘ��?g6����H)��іb�Sh�	���#G"d��H);��!��%��l�:Z>����t��Pך�w���0�����"��Z�}�ܳ����X"��G�!͚�I��]Ӹ��0��!�6"�oi�XcB�dk{ޥ���;�6�ϻ	O�ǝ��O�lnu����Xiʪ�2��^ v��<c��h8G�&�uC�L h�pj��@E�Z��~S��RÔl+3���	�mk�P�:K��Ʋ�G�|�:e�ɚ5*<^l�F'Q�����Y
jh��^�KՓ�����*�廵��L�o���:}Ҁ����Lv�9H�r@�o��s�s0P��l�����\��v���E`>�Uy('Ip�]XD�Lо���9�N���*�+��|u��h��F�4�:��^�48�8/}T������"��~��	���di�3���������(Y4q��bFeʈT  ۈ�)Z.ܕ֏逕Fh;[ �@�\�ߜ#mwK
���+�_p�9+V�b�$N
_�'I�f�}JzcUS}1�Š����������J���z��j�^"�����^٢g&Av�2t���K���3�B�d�̣5mL��,>��C�����%"�P�� ��|�|�q��+�؍�1�d���a�����x�	�,]��~�$���<	c��q�P�C-�V��<���\hh) D��(O�O����pэ�v޳��J��.�~����uՃs.�ދ�W$m��b'	�����.[�I�*�V��^��kds��}����ba���Y�Z&�a��h7��?�B�#?�Xp�=������3=9��/�Ѷ��]
�����[�~R�����֢{.�'pM����K�<10��d{��r#�ܱ_5�D *k�l��}gW�S�\�&t�h�]��NE��'�ч8�5<��-�}��7;M��:%@i�U�B�E�YH��;��p�R�g��` ��5{��xl�A�DA�?�iÑS�X�A�����F�/<f/�;��X��4����g|%-)�z��Rg-��3���y��W��>�t��ƼN�A�,�۱j�7Y����jP��&���l/c�4vq<�D�������?-�7�
��QZ�W `��ѵ�Ɩ���{���L����Ui�X��EU��>���Ta6V.sz�C��G8`S�"� ��gkLPv��=@H��MA����Jyp8�H��PI�N�bJؙ�.n���N�4��6g5/4���&��14�o��x�֊�T�GC��ė�
�f$EU�<�^\S�8ҨpKxڜY�)�)�'�-P.����ẘ'�+ ��E.����٫�,L�k�l\ ��<�1�,�hl��A$/��g��y��s��Tu���Jkm�tV��{��x(�s�rJ+����C��NxH�ca*2jy��pl�4��\��~lꊙvrPBu8��"����'Ya�|��v �/�BB[C��'��:<���]K�ZPod�r��i�q���S�%���|C�,	c
B�,�s���NݐoĦO���V�Y�d�f�H}N ��+��.h�2A�MyJ��n�QTPg&�)��b#���Kr��h�[��/$͊�^���(�;x�6<�X��զo����ׂ�����ȍDV�>u�"�������?���G��m?��_6���AW/���I� 0�w|7L8���r�W�T��E�X�s%��pX����X.�����a�쿲|jvOɅ�[Xj�μ�N���E
����Z���>��~��;�QpG�֧�U��y)�B����Xt`y��Fc,+��=N�psҳ��Ά��&Q�䥛�eáꍈ��7	������q7�J/��F�z�}o���W�n��ӆ�#GkkY�a��X`�V���)�y�=�bI���n��NTL�����bL��Y �	�e��F� ����r����ǻ��0Q�Y5���鏰�Ye���? �[&\yĒ/V�;�� ]�Z�u�y�$�tB	G�Ateg6D��b�)��3��)#i�
��#7m�;0��0�&��`Tv�
�\cI��6�S`��.�J�MT��1؀����-z4��1��g���.x��YPcK	I:BW�g8{1�J2R�+TG	�n���BlI�@v���G��������K�-�C��V�I��04��/�c%\���}4M׾� (�*�&��wc�ߴ�L�}��_�<t�s������<L��K���:[��7hY�z�N�i�	E_��n�@53�e�51�~�?>,��6E��'lS~>bͪ$��X�Ź�'ji��r�'b���������DaS���l�]�	�]�zW%��C7�:�X{)�\�[I����|:�����c���u�Ƶ�-�u�>?�j�-T��w/D�1j;�7�b��������19R��H/�����y���P�GN�-�O"#���!	P4��p1U�A_YA��\r�Yss�)�F��V��`��ww�;M�p@J=�B�����t�:�D�J.��[��UDj>^W~�B���v�@G��(#�>��)4`����xl�iCZR5�5&X.��5h�y��K��ion�bY|��k���/�Ѣ�b-ӝd���	��8)�K �Ț$I��@Ө3l���׉���cWP�$�@����{ʿd��ns�<x�!1Zm	^�3�D�r�T�
Խ��DC�:�����D�7jx��F,[hVK�׮��8/��d�J5|O���/�?r5���l�aƚ���w���|4����o�3UT�P_�M�k���$i����m~bF]����xf�d�'[�`�,.;w�8�mNQ�IM$��0r�[A���89�U�Ǖ�X鄦UI�Nw���;�7i\��9%�����b�4EZ)�P�?!6ԅ���c�9#~�ə?���/���1��
����m*u�0�+y4�P�x�c�&���:�KwZ���W��[�����t���l��6�>�A��7� �c�z^t���>����i��F�M�V�[�9O�(�욶"��`����* '��ő%�)���-~���E6<���T�(x�U��P4�r�������?N���2!/����=��h�#h��[�$�C��0�	��/��d���.V9���8� ���j�8h���,����8���Z-�� 0�6�^"]�h��� �J�IT��@�*�Vy�W��e��Z� #'j�$3M"/&9b����j�����X9(������&Q��T>���	1[ǄX���Mx��������#�V,�߇�E��ݣUl!f΂*Ng�+�M�W�II͹/����_� ���+�-���훕f�Pi�(�EgtvR�����7F�2�����0kgL2C���l��r<S���ފ���Uh��5!�+�v�B���qU31'oIZ��ׂ���
���4`^�M�~!.ޱC�s�&��=�D�2��󦺍�dj~`S�E�^�_s�~׉G�������YM�N*�V��g١�v��v�XJg�;o���]���Lߦ�.���·�9W�Ah�,'�1t���;_��_��z�> ے-1$���sV��&]�F�����6�ix�"�k�]��0nEA!����	,��e����tl�V��y���{�6�F�aV�盀��x�S::�L�^�qKIđW��?�5�N�,Y���[���Wt� ����w#^F���vͷ�P�Jq����E `�����N�Y�����W�3�ɘ���8�
g%v��b���t�������9�V��)P��~UܑR0f?�?L�=���_�f2��hH��<���~~\R�W�)hz>\|�ɫuL��K�+ �n�v�x��\�SMd�SS��>�Vh|��jv���ۏ��3R�Sϣ���-Ó8���>�u|E{��Sg⮫��k�.��>#��b�>-/9�������k��g`�t5�r�+��_+��=����!7R�ܚ�K��;�O[��U5���^�8�%�������hX�]���� ��4O58m_W�$��)qb��X�����Je�0�)&G40s�NY�_jQ�tp"���\�
	]�uq��:����U~V.�$�ps�=��I*��P�VlI:�וx�"4O����f�~e$�WY��"���z��qz�$3zʺ�)T��&S.-%�]�����C�(͡,�W�߰,����HL;�?�� ��v�'/�������!;i��Й�N�>�Y��!�8��*���EeP@��@�gZ	W9�¬g�2�����OQ�KL��-�z����J���odè��r��d�}[���qF��jGWL�w�OU�J����[}��h 4lHT4��v�_)�� ��|�]	<��.1�-1��pOҍ���M�����z��_�2V�Tf?>��a�C��N�Hd|V|؁��m;���N�]p�H��pf�j8�Z���MH���q�+�̔�,��l㠅�i�Ƞ����sd�Q�r�&Z�H�P��Ȟ�p���w�ǉ�S��2L�H����Y͠������Ӑ,�pY� ���a���t4��`�¶�b�M�$�d7F�UP/��׏WЉ@���5$���G4&ݲVK�>�z��W[��j����?)2�Nj�"A�� �(�Ҷ����k3YE�Pج�c��GAG�+��Wb�����SIS��f�v�[�l��C���{Ci�tpC*���`��T~-H���/��>ϐ('�<�$[���UX��f�r#���\K�8��|a\����E켁'j2�w</�K��J��p'ݭ�JqNt��Ȁ�ٲ��̘W�5v&�A���7�Ǒ�C�^��}�N0΄{n�"��B\\/ٝG+���^�uA��I�m=���_�5��e� ��V�Sr�_W7c�3_WiT1�X�GϿ<�,Iے`�nIU^�w���&N���f����!ME��~ʈyO�
�ʈ1'��K�f{�%�D���s�g���U?��K��i[��Y�9
^o�f�������C��Fs�$+���?����^��}�3&NB����Ј�)�����{�Y�ap~�DY����^��cp����u�����]�~�'� �t4@g�����V�A'.]K�8���Rsa���&�h�rPf;w���f��)ҫ0ߦ4bI�WԉN����4oRr�.�@�ʼm��[y%!� B����%;!���K������3�`�
����{ְ�<��L�0Jpڅ�cB�K�J�d�L�_oW�(��K�2\�r���R]�L�%g4����[�uh���ũ7{�T�X���<���׊�Y�z'����}�w�Z�Vt�����DY��^T	�I�LHR�F���b�QT�T�a�~��e��WU�.�"F?�ХC�]���4�����C���r�-���ȩG�w��M��y֝t�-Z:#+��d��||<�I��x��e4f�
������m��5����t}5LU|�vY'�ߍ��rVA�%����5�l�E=X4E��-�2+Jw *����V�2�U⚲�ĳi���zH5�*�2�� ���G�@���0�,`�M�b��q73������O�n�����,��ǆ���ڢ+*�#`B�Ò�Sx~]�(a9v�:h�3x^���Cbs,�RV���X��9��aj�ѧ�(�~�#���۔�LG�%�L8]����)D"���/�m�,�z�ӓlUh�]���MX��L��~�u]�0vA����W������u�O�&��;�hsF7d֙ �6s��Dm�ӟt�S�����lt�!�&���e��'F]���]?Jn 7���U��
���/��M:m�+�D��{eǭ�H�T
�'�x06Q��I.�;���} @�c/h��1���1���+� 0��(����;$�ۻ�ΪM��^�����$wLf���ƩM/)����'����תB���aܪ���?S�b�P�&���]ѝ��>��U��I�3CSi������9�&�ʍl���%����$��h-K��sY�u"'��dͅ"�O��ǅ_$:���<�'4�o1�k;v�x$�V�֖Hx�Bd���Ï��m�u�2B�|��D���r�(f�2?F��h(��p��}�$�a�k?Jo� @�N�1��	��YgUh�� �0IE0j�z:`���c+�����ETR>�jTۅ�s������y�Em���Zu,XL$��P��xj�I�:�51G��h�,ů�!a5�fA���A�D�D�)��8�BW3���%9Y���������c��rM�f�N�/0i)�WKϬ��Y�t'�m�����B�,`�{�����R���%E�ह�Y����t a�I�{��|�Ȧ>�b2�u�������IV�п`��,2��Q��;�wE�1��'���m��g4w�O��:���Ufx�Gw��j�o_���?4��+i�ީ�*0_P&�j�3�iK�E9i�_�響7Z?.J��J�m:B�c�
�M��	�L`@��L��&_���K;w�	K�Q>�k�T��1˙
�]��)�;�)Vo{��m��lB���$c��Q��N�E�<����U+�|98��E41-�E+>����D���c�>#3��b�i�T��W��V������<K��H��~��9{�B�ѹ1�K���4�8��]���ՀBVi&S	G��N�����A�Y�}� �hL��B��i���k�~���/�πkv#���%��qT��z������I_��^Ƕ��5�s���v��X���@�����sutوs��q���O?+*�}������#;;s��"H���� �|�@���RԒ�'a�����9	���lQ�H��s�]�͂��l.=1W�vQ��*���d�{y�	
T�a�ꕸ:^�yp���I5��\���o�"^x�_��Ӎu�?3'�X��F0a@Ѱ�/0�o�_En��K5���T��r�-�od����(�L�4R�d[�h8�Т�N�-0�F�lY�3q���U��O�X��ޘ���)B���X�b'L����`('��7�-ۙ ��O�4���V��.#�I�6�yh�okm��O�fN���L�GF�j�/J�9}_�6�\C,�wl�9,��7�����}�3DK����޺� ^ڧ����?fv�P�l�c���k�E�,�w�?�^��v�I'[�m4���b-��$�2���Ѝ���E_��7NRx%��&�+�ˤ���Wڲ(�?L��g�$��5�"bV"�u���;����wh�%L1��'�穫��+R^��(�<�y�c�ݸ����>ۋ�x�ܭ(
��Z<c9����y!Lg�ꎡ��1j�������}��M��֬x5��}&�����C��f		��r��b��Z�~��eR����X�k�]�����bPun&�E�J�D!qu�����iZ6�Q�ʅ6m�*Q3|s�^n
)��L+[�_�����=t�5|��<h(,�NM`�2py�)L��q"���L`�������s�㄄Qg�1x ��8 �qg\�&��c�oC)c==����%怘��3x���Os^��/�L�#V��{�;��ak������Ld�v?S�,�ɣ]����Y�M�')�����W�$@\�<��Hc� D6H�/B��t
r�'�IB3؜,|Ȝ��F[v� ՛<Ey���[�2+Ā��o��H��f,�䉍���� ��!6n�W�Ck�6ӿ���R�, F��2aW��\�8-�����,l��/N%��XDӒ�0)������DC��������,&�%;���8�%ՍUi��fU��#���~с<[������69P�5o�q�G�J�/�h3˅n��HRɊ�7h_~D�C�Rv����mm�{`������#�{����F�7<M��p�V�9�NW��xu� ��-����b
��x(��U�&��Y!�S1-�.�Ǯ����":��/C�i�D�*�E�{��=��7�i"+GVU�|Vq �ɲ�� ���3(p�07��U���uE`�V0 \N/_''"E:"OW�ZK�f+=���}c��8~,��n`[���7hn�����O*|ۄڼg��<od�WH��z�r��aa=[s(!q6�����j����M-��y�@l��d��@H��k�M���F�-�#����	@�L���?呟<��! dxaa;���D�`���<�n��ۖ��mP��P�x1T�!��LK�B!c&��-z�Ա�-- j?�P�I\15
v�p?:`'�Y�́����L�o�)�=M��0�2O/?.*��q,�ȩ3�@�[Z>Y�0U!��+GrU���Io�*����"�t^��Ŝ�^3���k���a�Ԕ��Ʋ8%�|����������鬅˚جw��7���pr�+��{����O���;�W\�/V��τ��z3��x3� �7n��B��{�K����,���EB�'T,����-a&8��LAG�$C�CLB�� ��Sё�'�X�kQ�VvA)*���̳���8Z� ��fv�Pӵ�+ր�b���(S�S��	�E����XRr�ǗDv��v]4fKR� {�U�$/�fR��}hӽ:�EA�,���(ӌ�̸�	�#½ڨ:W��$84�8�w��+���Y���R�����a��x���V&V�0.%'�ӆ�����RUx��&�G�W�%����}�<�`����?}J�����,Y��y�oR��]�~�;7`G�����[d�U��U�b4HI��0�E�T�r�K�ȧ�+�c|-`�:� 8w>�.���vsт%?���9/U�}�2\2����Z
���y�:�9i�Vd����	�x���fz��ބ�I�6��N�ǩ���71�fj��=�����ZN���*R 	�4�Ie�)�0����+�����&���欯�+,�ɜ�"�Te&�_��'}l�\�t�Zw.�񅀎k�*��ěpǺ�7Y
�p�ݐ�d�~}W�<� ���5�>U*�8<��M8b��OB� fF��nm�ή��mN *d��3l�Ⰽ���{�2��a,��Լ5���p
]��v�~B�}���y�:�Si-v7���_����s�0s�6`p��"�oz�r%�#-�;�m4�7��40�G9Z����TI���H/���?OW3n���q�{�=�(2�`_u���.�M�G�N�(���噣��B&/	�շd�+ ٗ9���Rg�~�w�)CVNd�)� �M�L�Zx�Ɉ�:(!��g4[�=�"_k�i}l<�(�T׶ae��_�<O�L@ϰ�v\x�4�<��j%��^`%A`�d��H���b�y�H���:�z�wR�!��:�K��V�y���p��k"0���b6d���R�o"h�!M.�/PV��h�jfr��^ǭ�@^�G+�>_�E���~�_��U�#8�>ԋ��f��������D6�������6Ю��yJ8Z�9�#|�4�\l��a��.;�������ãY�����5�Y�<څ���oJ&c���@'%je�9��%�\��Q�Y�֜����b��x���)!ls�z�)Ï�YC&��%]~J�����e�׹A�^�^Wh!����@)�7U�W���:��翨�	J�����C�´�W�Q��.�B_�D��	��� �S����t�JƜ8��1I]�X��-3�x�R���-K��]���76��>�2[X>rOuڹq����LW�M�^����^{xKR��7�#��r��7�}T�:��f�j��&���	:�7e��2L��~԰�/����T��/C�,ҥ}�%.s�s�9tC5b :
��fq�Ou���A&Y`l�l
9	p�I�wN�h8�P�q@�@ts�9.�F�fc�t��ع�w�+��Ϯ�ÝP���m����Sن�R��٥��w�e��dK,-X����=P�[�=;�ŰQ���-�-b=��q��%{�@l��
�������i�\���V	]{��?g�	�4���sU\D1�*]h�v�X��5!�Y$$�E��۵]���(Ä�	W"I�b"�՝�b�o"�Z����J��c���a�8
�M��"�u���8�
� >�,&TAD�C���ˬ$�"#��{ױv>pR�_��I���(�)�� i~DU�5�9��,�B�$�0.m�J5��o̈|8R�%��a���J�P �gJ�1����n�Ǭb�zVQ�W���h���֙�:����F��+�o���Y�T)[���ґF��y�n?w��j^����{�.J�ߺ!Z��*s�0V���f�ݎ��}���v�Gh*�Q�2?���� ���Y���H������y%����B�����n�4��.y-(%�dM�i��FuҔ���Q{`/���<���J������"��LTe���^��mY"���n�iv�!;-��%F@mb��_W^������ȩx]�Ye[aE�:�]������Sf�9�M���U�pME�r ���ŉ"�'�5�ol��${��X��(�>9L_'�NZ
:��=�S4��J���RZ�t77FU'�!��r���.[�gЕeo����֗q��7��}�%�{�%+�V\�������Uغ���w�9X��w)�`��AD$0��8xX�$zq�����7���;�d��A����-�Ex�0�Y=!a�+��j�[��ޗp�7j������loֳ�,}lY��j�����z��˜��zq�h <Y��30a�RQ���bF���sލ�aG*�}DT��;ƶ,6���:9�_�׃6IG�����OՁ����U���Y׾�ʩ�𘀠a�����x�����b�ǟ�B�w��Z��1�_]�T���H�@�����Bķa�n�Z<��L�7���i���������J�3s�-�W ��y
�lT&!v$?�>3�,h���3Y��&9wY��q�<�	�4 R��j��Ŧ V._�JV@��) ��Pz�ȞnMS��n|�W�/V�%�Fs�,��-
Q��+x����\�S/�^zT~jd��nk�{2��8����](򾄵.�ׇ-�I1��~�ha�ë�e&�!":�()��׮��JE-l�VaQȥ�e���"�U�o��vY��7�	0}�6��k�&�	�?EAV������o���\�K���֕�0�$&S'�r��?�s_ڭ7�}�10���{��`� �8k�~<�+x�����yk7KP�X5����ihk�a?O��)��V~�A��$�z	M~��S����bk��hI �tl��,N��fӋf�� !�M{Vӝb�!��M[�%���!�HL�?�~�&���+F���������ꮛj�m�L��#)Q���b�$���٠'�W����\��yf�KH;�yV�9�D1 y-�������}�:̴�yw;�/�Mn�
���u;�4m��	%��sư3����M�}L��*mIʈp<���+���:Ides���=��o-s=��0����bG��|��$NB�<һ���֜˂`���qq_t2�F�-�-W�o�+9��`����.�na_����W4Q�p:^�ҩ:�Ĭ���z��ڧe�o��B��7���p����_��p�PM6��Z�6Y[��o~j���?���D����uY�l��w����w��M��Umi�𜉉
��qR!'t���R�pX{��m�nv��6��K�7�pl�QD����W��2Q��g��-�3ł �^E�5-�O1���F,�~U�E�;������=i�>�2*�����q��A4�B��$`��VȎ����[��au�	��(����j~��?���҅s��F�	���<8F���Z�Vqb�Sd���ϟT�5`sx�	�qR^�KKgU�2�eǕ���U��U`��SQ0g_(.T��je�����Ͼ�EȻ0��1_~�@V���%fhj�υ42���]䅕�M7�fx�H��3Vk��D���2H��� �Xw�x�\A��Y��Q�X� �^�e��.�� m.l�Us�ST�h�P��d8#�"+`K?���m֩a��g#OҾ��EٽȈ a��ۀw�����AA:|$������V�Js�Z�Eirm�r��'7,�M���9}�οMo�5��.�#���Z�����lQNO:V$���0&������>�'�8m�qt�A�>YQ�;��I[�2�w�Ϯʠ���a�) dN�E2�����l +n�vPͲ��BC�Y�RD�L�y^F�6��e��ֿ�g�H�ʤ��p���w���,���?���ZB�ׯ2����G�<�����׹�Cep�T�ϕ���S�(�鿜Uj�Ң��"Ыe�Ǌ�L���g��5���҃I����+��n��+b�0����4@��%
Jp�IL��d��/A�|��U��/&�2�؂#P��y,D�N%l ��s.�s�����1����su���S���$���X53,�)�~��e����p�����=k���x�T�Eꮩ� Y2K�].T���O��[E���c
\6%�G�ذ'�R���Ř��eXn�Dr��^�-�Ũ�I��o��Ԏ�#�OLH|YL�	�M/7'���۽�i�>���sN�hӾ���0���nr�d)|��Gx4�������8l��P���s���u��"���R��=4�"c�qBJ[�w|+&��.�`�3SG
U:�3fn'�/�����C����q��< �P���DP'7�����O�$��ȍ?�����u�׍�&.���]�:D�+��x��~�g^H3e���r��~P:JZ�My���1fyV-�:k��Ӓ�hf5��I�2�O�?���	�k���J@��W-���HB���P9tM��EG\ٞjz>aO��}-�9��OĀ���i�%DH��j�欙]�H΁S�4�����n��*�������?x�TG�����+g�<sS������S��>�1$C����<g|^z�xT���Y��\x`ǡ_�Uw4k�F�3�:[�����0�jގ3�CAiĎ�4[�����;
AЙ+�Y; �	�%�
R���g*d��q:;���}J�n�*�XFCaJ$x����I�Q��OT^��|B�ZX�)T'�EPr����������ii�>�.AO���ؔ5�|���+^�gAf��B��[�yN��J�.�rƔ��r/�)��%A�U�
�[�͜7�"2S����}��}@ީ�s7�0�ba��w�����p�����_���=�yd��˃�N_(�Bp�5�GW�1��Gm� �NL���c�M
Q��/B��QBl+�1%��Rد�|3?�g�^�1�lv��R8K4��@:�����9ё�)�Ѳ��M%�lK ����h�-�W��9<�3��32��u�s��<T��a��6�.)��(��k��X�}3����
��pc$|�Q�������[c��V�1���&����vjH_�v��rܻ�C��I8����f@�q��AR�]�?2	�kھ\���U[H7��_�A
0���d���v�����X�&z����8�3+��c��u����5�R�� �<ڤk��lں�c�ڌ��V���T:��JyG�<�]Ўao��u��)��g�^�u�����N�FP3g�<��3-�fD��?2-�b4WakF޼�8T,4��HR��3 /���A��5�Y,k���Qs4ef�K�q�}�ћ��A��MK֑R۟,y*9�PS�$P�l�>�K�b�ߡ,�^WQ�E8F�3#�}*�� ��1L�~�A�8�3�ԏ\+�i�l]�a-KTkp@_�*JzGQ�AL3�\��{�W��(y�#9�ʏ��̱l�}��/I��N5 `ӈ]��g�箟��C�C��n�U%5h��cIK��HO W_.�v�jD�^l��EE�Ubۏ��2:����0�4��H��ǭiu�8M!�j:��`��g*q0KႨ�{J����m��C�7k���U��2�c�j��S�py���k��ܫ[T�^R��w0
=>�V�x^I���9�d��� �[@�MC$t�#��S?�~b�1F��d)D�OL�b�N��jv�q��O2uO"e?��ra,^ ���o�lШ�WMڮxX�o�	׭�� 3�gC����Y�������F��R��]�.�7fE���}�L�[�3�IrD�d�x%lR6���~��#P��� �Q����
I�jX�3��0�!���$ݗ�z��`�t��#�R�+����nӚ���)���3�3o�;���]��s�ft��2�����43F�[@�[ ��2�b�t/0��H)��d�r��Xmm<Y��4Z)�'O�4<�����69�����W�!'�G�����	��w���2�	��=���ĕ���T���l�j7]{q� �b71��]��G&��Z��	>�0Ӓ<�ǡP���^����v,���q���0�X����>6)��4#�`;pRt�����À:�kgKt�G�l�C ���\�ښ�V8�<���
%�O�3V�,����Iyd���[�I��B�q�E =���Q����K��d�,�v����r��u�k�Q1��@�]	r��;�[��r�j1?jU�4��S�̠�1*�pF;�9(yU����
��0[�Li��!Or"F᩾���8���Pynd ��u����*�A�N	�����0��>L4\�o�y���#o��x
�]!BYk@*Mf�E]��j�&�dZ���9��8^:����,�]J@N���wJR6�����=�BnV���T<�Qq�|s����\g��&����`�z�G�QZ�n���0?�Lj���xv �IPV�%w~��ld�v��t{i;���n �����K�V��i�]�쵓�T�����X#1�����\#��1�9�~��>�J�MO�ζ8w����?Ѭ�v�Ī&t���Myvt���3�!��Ϟ�"�b�k+�h8�1�Ki��������l���!�}z��-� 3�0G�X�2�l�}���B�4��d��mf
�2�?@�މ'�*H�=&�j�S�gjkBU�������o[�� �̇��J�j.�)�&����
C�����ڭiqM��ļ���hV�N#�g C-CR����Qnbb1N����4��L䖿RH���H*� �7#>y̕�+�;��./ɧ��4'����j�h`�s�#=�I}®��.mr#Z�4��uw����F�A��O6\�ssQ5H���������`Tg�V�H*I6�i;�;徺��
���c��]�G�*�1Χ#���8�kh��gc��PppH���+��:,B0.g�)!���v�ZV!=B�U8���ݰ� �mA&�{g�F�>�l!� {/VZ�ȸ���+��j����C䃣��28�����r��)� /O�,N�ݝg����́�+<�H�&��ɨY�7A�&S� ��_�L�o&�LCVv`7�[��B�r�턙_Vy/����|��$S�6E�5�u�+��]��@�#���zB�h������U�&��:��)���P�i*���4���r`	�<�&�W�5�m�|.>�Sۼ��
[��w�d���V�\jYz�R
�i濫�I�zl�ϯC{�&�	�sx��o�`2��Rd8I��U>H�3�zw���o�_+|X�Q�S������8�P�kb�FՀ�T�-o@�gK̙�|=�d��W�J�p�/ZG�!��[���V����kY�1]���������w*��"��E�,z��n�
i6w���3sHShˇ�=m��WU��w��0�4k��~1_4���q�h>���' ���hp�7����0aafT�!�,�卪�������e;?��5<fЛU�t��N�7Pγf�f�X�m��'�v���U2cu�(
b�D�M�,�8�0�!�%sxc��s�d7��D��TJ� T5��|
���	g�����Q�zc�
3 �3	�2! JT�0�	0��	}���(��������!iL�.��	�� �ɟ�mE�RZc͘�)�SǦ��v'�s�	���}��$;��;YΠ^YĹ�h��>>P@֛D.~=�ۄJ���S����%/W�9�Y�b�_�΃"o���ڨ��~	rblj��gShU�à�@�{T�_��U[���cm]k�i9뻸�0�2�Ӗ~(��7g���.o�&��`��$D3�a-�S�;�+⭊ӸX�A�-�op�Xb5�7�IǴys��.���Y��|��֏9�l�'�]2~��F�I���Ź;�N�#L�0v�f%���T���5�.��j�?ʑtM���OG��-�2��(�=� ���qZO=c�`� ��ΰX/gk��&s'�΍"��;�?nv%&*�`E�
hH�W D��> '�`�5���ӾyH��<�Of�q:qZ�#PC��t�~[	}a�6p��v�� \ �V��,���]1"BU]՛����35h^�P��uqI*���?<'�;^��듑�iAgH'��d�o�#���7&-�%'�n.�9�ݑS����3Mo�N�C��PiOE�#�҆ejZ�����!��V�OkEb� �9�����k�ѐD��0��Y��?�j�vK%x0�T�+�da�nOtd�~�J
aɏc!�P���[���N��\r�gKA��ɬ0Ca5��<ڦp��(��%�<$��N�a�@�Ӈ����%��i7�<�i3gE�
��w�&�e�䢻,��"��'!=�|�W7��t(k���c�C���F�����咓����̺F��F(���8�q��@��n�t-��e߇�[�K�A~ug}��$��T�D�e�wo@>���`8	(l��qh��D}jU��0n����|�����Ԥ� �}��Dm���.`�G���fl�`<�-�S����>�嶵s#s��VƧ�:	#��?V��ᳬ�V:�]$j�HSň����l��0��;���Z�t� s�� V����%���0����|�b�L�"�I�Mpd&1˂�5�_�qU����U��n.����n߲sjݵ�(.QLJ�E�l$� 
>v���ֈ���Iو��Q��h$� q��gͭB�iHu��p�z�-�� ��v�+��>'���bv����0�j���GyC�[:W9�綊��f�-�Y3g/Gc�5��	d��33�"��K�;s��Vj�Z�� ��j��όh�#���ؑIN��!��,�>kc<��r�4�vZ,W��S`N$��"J}��T�9�*��A��t}�@���U�ԞB호��(�$�ojGS:�E�F4�!����f��7�C��?��ܟ��x(A��F5h_���w�.
�X�9������MD�&&L�=wo�MVFݔ���������nN���NL��3	T��Ų����l)Oʒ�j]��ov�@F-����'���#��=�&S���]:��C�\A	)��ʨS6d��|�{��fC�>��I�*z^}�,�_7�A>u�ꝴ�@�f3�D�F�ung���;L�Ѽ�-�z0P��f[�P��!*58��������dxq�������sz6;*�i[�������J �[�ҍ��v2��(�_��W�U�1G����G�^0!�"��u[�wx�ɇ�(U�ع�E_�Ax�z����5u8(b����6��3\�A�t�[o��R7kl@���H�S*lEMY4λ�m��>�_�c������r�[\y��O��Cn���<���Q$P�qp��T*d�Є��H4���ӦB}���u-��bG��=�C�O��`��G�����(з����a?���Ν+�^d�i����4r�����G��	��Z��G�]�,Gj���[��G���o���N1n��$��!���8L�lV5!w��P��e���Dq5̰G��Y�X=��h{��QjwHaE
j͝���JM��Ӓt�/p���"�2�A��oZِ��IZF~��������8��S��r��e��[��t�X\�
gFP�Z�)�kv�ڵg��G�d�Q��:]�#4&L_���	Mg�z<�6=◉C[�3��na�N���$@7.�W�dV(�h��QELɷ�5�)׬5৏ᔣ�=���!���P�1�B�̿���е���X��4W��1��	�G��N9�n�?�}�qQܷMR�[��+�[�d7,M�*x,q.�3