��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,h���~�G��G�j�V,=�ԸL7���[��"���:mL�Nn6?��.Vts��$U�S�C��I�i�j�붃�}즊�üå%����6W�	����:�-�=>:s����u
�I��3�G��U��Q�����I��F���bHiM�x7�$c9�ת�cI��h���5rTTg-�z��;5�CkB��f��z=^#H�`v	���R;&[B�j�Ej7�� ��j�GP~�Yc��nQP�*�_r��cE�^���&կ�Ҭ[�'��H�����c�P� ��F+�PQz�<%ٯ�(QZ,�n��2�{�a�\�!�vI��z�:c_9"
�6<���u�|#��	�nt}��){��ދ�y,���h��c,�]�� ��Dæ�C����jK]�`сP!����1��e��7�mC�9��60��[�Vj�O�'d�p�ݮmΎb&(�"�*� ���B݁�ik���09v0�3�p��-��$rq�lN�[�ƪ�e�ɮ�����^X��l���/s����u�D�aQi~�1(wTYF��P>���E~�=S{w���耩z�F%4J03����%�X��&ۗ3�e��ыo_��Fl�m�N6�����'�Q�'�G�����\-�qR5������vx�݌�S�H��Y?�{nW:ђV��S@��K�$	�����ƙ��y�1S��� )�7�`o����XT4;��-�����!�U@�N�O�OuZJLQ�Z�O["����j�R�bu�a��V�|8� ���6��g�`i��+)δ�]��`�"0��"(��G+*��2�����b�)c��y��$��Ǖ���Y�=����Q�T��V�Qg�o�H�h@��
�4$Y6Dºֵ�=��P���py2�P��*pI�֩q��5�хڼ�]:J����A���5��3 �z��fr��Dɫ $YK�������m�];�,�u'� �p�ݛh��|����+���Iq|��5`���&G�Z�-L`��=OZ��N�?��؆J SlC����OI�%(�ޅ�"�[p��R�x�3���?u�@r�
6��W{Let[ ��bY����9L����1��� j:���ݪ	8y�������1������j���$��쪥mr���/�E��O�:k{r>��̢\p<�f}Jϩې6Xc4Z,p/���p����5����*&J+ ��%"Y����@��"f=i��fEǠ�K��ߋ
��_�`�5:�Hٝ����[�]`�W��{t?�����C�O�zǷ��A�=�3X�:�&�cS؜��W?��d,F	��y0�=��q5�Q�a�ڈ�#�������y�F��*�^`Ԉ�Z`���I׋���2�BsE�F��|M,1�]g�k�W���Uȇ�
�d��~Ѡ�|<gbQ%�I��|�2;K�������G/�5�|N�X�Q3*8�/`;��#%ݼBsV2b�*@]!Y4���-b}�0o09$A�qp�	�TQ#��m��z;�@�*�$(Kl6,��b�!��pw�%��"�DT�LS��X0Z���Bɗ��N!����*��^^^v���!`�)�D�x�b��i�;�r���ݡ��ܣ�tO��!wkRP���Ҭ
J'|��.sT���#� V!�����w�s��M�(�S2!��S4�$j���xQ��͉���7�&��`��f�Z�TT�@������O�-��H=�E�5��W�q���t��B�`�n����'�2��5�~{LsF&J�RQ�{v�8���Rm�|�ґC�������b�F'l�跧��!2
2��G��9������J� ���$��]�7�xq�/`��Ҕ3�������ci)��oE>�V*ܸ[�2Ƒ�^2�ˬf�o{�:�*��<B�ҔP��������n(�Eg�u%���t��Opuر�H�9�d}υD ��Mքf�7'�(ƨ����8y�V�����C�����&�8�SA]��Xl�u�O4��d��ڿ�-Y���Pu��ߖ�E�)e�]�zb4��-XH�Ҕ���n�+��(�?�.-sr&�K�W�����3܆l
p��PCg�3�<-�/����vdB�)�H;�|��(�n���X>TI\Աf	 s�"v��6�3U{í�<$~s�[Gm=�7Eyb���`��񆎣M�ʩgt7{��V'B~͊��O̅�������>?hc��d���D9��ǘ3��
�"�����wJ�=Mu��`#�M�r�}V�6�*�p�V�ZT���#c��y��kU{���G?ɶ�1J�9�$"��(��MW)��o"�i׎��r�8��/P�鍀	�Y�J���[�S�,��j��Lʄ(S/��R��+�(���h�F�ɚ�q�HT� 	�)���m���꒙��o�(�o
�X1�M ��`��Q�	Z����P����I��M03Ab�/����\���^��ъ"���6�4f]����0B�S��GQa�j��~�OY�1j�Њʔ�~{�:Tt�]Q��&h	j�WZ��EA�n��7��	�08"A�ĖV�*��vo?��?\���Ɨ�@�㕛}y�%�#F���q��]�E6)��C�8��}��^��s��i�|��9-��G�aU�}��+��7h�#+���B[id�Iz�3�i�6/`0���U5=�/��<�~�/6�:�A�vJ}�܀���J�q64���sM�sUH�1���k��{�6��i{]ad��L�� AWǬ�cm�iL.��Eae���Zh'Nn������f��7(� 亶Q��Y��1#;tC�hi|i"�y�mЈN���w�2,�����O=·�/��G_�0Z+<�}|�h`��$ ]�c�Y_��B=a���p�|���`�C�u��5�&e��4��8�Ά�cU}����>��W-\-+X���D�ff����lY����%�tth�K�|Qz�i5�k���&ׇ�|7���G}��EYs��4��B<�d+�QL�S\B�u%�3 (lV��O46_���rk�y� 
����tf��)����](��ؠY�g���ɵX�8eX�)i\�ېy���[r
/����(N����c�W��x�37�3U��5��G��.�;�U8���d������8�K�`�8ڔr�yl	u�5�!�cx!���� �p�*���E*ɀq��}Q�C1b��E��6V蹐@f*�F�5&�$$�`	|&K�$͌6���24��ւ���3�`�]$�L�o�