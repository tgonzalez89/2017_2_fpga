-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
EcM7784d/fVPOpHKJLUl5dsyCtj6qWc0obAJ0uUj/UbYGqOF6dcC2wab74vRxMeCG/NaeyqnT13j
V3buKhmyZhaYJog+808mmyTNWwgnqlRxl6rrda6VI5MZsjaQHp/ExaJPWjxzaRAOsHFo0/oCNfCk
Rw8g5C+5KE5v2J0Jz6zI0X/0edi4haF30rgooeGB1GpLGE0Zmr3+ZLkHBkc6LM2enNFsKPry7B+U
H5AxnXVlK1GZXzzaDcac3gnZ+GxukJvKItp7V+sWikJVIcO1aqj3t55WmxKPqayS3geWLRwv0HXP
bjKs1/F2gyLO+GCMeVadMsmdYvWhB/O8zNQI3w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 28752)
`protect data_block
y4rRBGpUAHR72lDcs3NzufpM8YYhR4jSWl/igUjapU/4Vm6FJy5q74fioFDvBusRjOqbhrAQvCdA
8rSLYaH5bRRyM9za105+FaT0mLb2UJqG2kQb45VGKq+l4LKAOM8uIqM/fh2/2xNsvCrBVYJhFg7N
2Zi5yXQVCbj95BdeotB4r3RS6WyrPIZkkzt3tQlzyD+HSeNo+jVSO097vOS4PS0JJ+LaHVCpgtEn
0yXpYc/9q+ZTF1i6EdpdQAClSEdwzJjwKe9y475CRe3wI8vIYkPzTNEVBKZ+pKTMWPoi4B5NO5GI
N6YuswO6n08VLVU08+X5TdLmWNOWrM2N3A4no7JEfqfLtryL3w3p/kNrZ+uPs1aaV0yq6xAIXiWE
yvj24eMBVnJm3WdAmU7KiUjch4tYeB9sW/3KIF6tq0ojQLrvlDZL49k62lB5UBC2pXS145Eu3R4Q
zKjfNG1ei/8WXz03/GrBXO2Tmn8qBKFwwdrkmF0eTubfvkbcwo262UDoKAoGLc8FuGWjXuWqrv1q
eP82bFI869bO+pbNzHr5DkirATN5Gy7OdEqpRLiW14y8+OMzda3wxsv2Xk77hCkm1htLo21THdh1
5NbHQAIrrj6vDqOboQhX1bk0ghvSd3+Ny0ARuWui6Vy1zmh7sIbWztx86IYiJNHPBkNiXuv81DJI
8lfPjk/uOl65vzp8yQJFTN2ug0K71i0Bx0SzJa66mbBQSMqVtNGr10eCOOUtnXfnSjtU39L6xs6Z
jCMPBMGXdcDeIvjtkfnnq9wjs7sLix/iAJmktBSIE2wBw8RPsqx3MT50UIEyhDZQoP000uhP4pVW
NPUj4nNdR5w4Dfcb15l7em9sAzy3i5ZlawDI9ioiso54zefalfTWdODsLVIjN/1ru7bn6pPc6udD
fb/UuCCAwGeKh7PmZ9+VkeeB3Ov+gLFTEmAj3VE2dkk4cL+G/5SXfzZIb7kuKfU8rHIzQMatGyCO
gi953Tq/anMpvumXS3k0r8iHs8syZ1syFytPNh3lEzjdDtgyBpg6S4d3rGMVzmprMMmKjfef8YKJ
6cUIrWHwqKQBouRXQSzB04i3IOwKJRRo/u1OAe7b48EA2ygcKmup0TCw9KuggVmc+Mrzcknz9D+F
BggbBuEFB8lDPInF/pXQzmKQxsm9YgOELBqxC1JgdzbhXcjmsBlK+P2CIR6u2tU+WIi41fr9Vf6H
bFgxc05c7mYHFgtKaO+UCST6gF0KFcSCBOPQvI5rsJmV85JZPAMOV/uH53Lq1W+d9VVvqwtj82+D
6mC72Ew7SBhr/MIGcRS1h1sRsViTWSDWMaAiCgMRQYnrt7c7cfgI9pxvh4EnRi/OnQ2y98Cq5es2
XErixkJsvoal6l4vZBnabRhsFQZxc6lUJc8SFNbhpegjElMTAj6vYaUjohfI8s+OqMmTyF8tvrfT
CPwLufqIJrJuo1p0rdZr7W4t54SzATOYItUMMTST+GEIA1btcSd/DrSZcZTj1b/PpPe+D+Y/RCbg
V6Il0htLgbmbeOmGAk96Cetp+z8VY1f9kpFyi2nsQr2zupaGXr2fX7kOIOwp9O98/Y4WYw4w6i7K
LJgfDjbpSazhihS+cdIEJzbFVRNzwfkTZ5zFqKClEcZu1HPzOxhUNCPLRLK65EPPaZFtNp/NViML
wuZVcWkEQUSQZPSG8I8L2uHmZgmoBuJpUyX8e0Zj/oQNh0/yt1mGfoL35Vi3TaUhUF1yTk7W2f1M
ztK9I/lF8K5OWrFSRdJAkCnhOB1M6aCoBKY0dqb0dpjYU5HAG6GVGmKZlki7UFhPa7iW3n4rmtPW
ToCU803Uk0+qB0lFsAj2DcHkB7tRoCTvNsPWmbmQUXmR4++aHrwRBUmG0uyV699PQive7GeqFU1r
d16Ejs8fTFszkdBVNjNA9iAbo/Ym8VHwHxl0a2MZv8Jc18AlSF0t/i+oGRypiqXSNiP3o7W4WqkV
WIYH2HAcfkUaS03A08eVabKf5SOjaljmFtZyCzon1/KAf6Pbz3Ko+UsVq9rzdGM4nGMbvm+vLLzd
jHZOQus3qf1kxqDqb/sLsm2nQyuA3ZOd4mALm+p4l5ZgHJ/apbG0k13zLZ0qKhEyTNkxnX2V9GxL
NIjWtpyM4SCbHkyjE7i6dhdsiyNDv9lC8ZgNXliW9hc0H5e5nhVfzaxMFkrB2DeeFdKWlgFyQgEl
sBu+G4IGxpvbIRorS8+Nm3Af9wB4QWvnzKLyOnaSRjCRo7G8xdcMHX2MREcLWtoS+B+XonEfxonG
PYQY45jdOvsqVfkQlG8qVjIuochf8RqCNzBE+vL0Q7rE3oYbBLJzLBRfWN8mkYJJNRINxfndT8nv
ArU0SEeXKJRzK2m2+123cn+lLtWYMQD197a2bRrXNEPa1oGppql8JsYBSL4Ny4Tz7NaH4sS4Hhru
IFq3YbxJ95T1y7q2SGw3DALjcXPC41mQbrP9NV3pw7WpqSuIzDfwDFFWfprMQLLK1ddUB7dZGzea
WUdMwFr0ga4pekO1gsk7E+n6e0vzuWKVdito3FjYgnDKEAC9CVjvZTEA90fbXr7aGl8GRRUyETbx
Z/7gwlmQ7uPd/+fBMmQ9W1YA6cXPK6CQN6rn/AVNQY1P6936eaX7aTESmkaWIEzj3pS/V8DY5yFS
pycpS0+r8hiJbMoYqJjjDbhBQ/aORg9geIWqdwLS2pzrEAM6pxlwXWRnbowCwsepmj6WU3zvjYi/
RCpm4isDKlgqSMlC6xwta+um7ltkiorEsTySsgk579U/74DjR4ntR6+UEul3bA42aW1niiT2DqqV
x3lF1m62kFQ/35yW9uC16ddsUTR0GbsO4AbnFXzeQ0aPjmMpBONyML1eGJ5JfGvXDYUw+zSl2HCQ
zx3rJYPiG5CWQCN6Bghws7AhKqcu548GQwiYVgm2tVcUwt7/+mOEajU07+YrwYOu8QRpTRTF3N3E
wz7/rCcXLBmhHES1AGulgjoCMZyXCPMezfXQoa2oDlHS5lXrrNn4KR7hSHnzXQ0D3APSouqMfRH8
pHWi8D4ILAweCtzed7GhaY3CqqCjJRNAHqc0npOU05RqDFJ4EgyXkropQYAhZlizCjQ5MGOex7St
lbQlHqHTGOOeKSADCYFdwnd1Q61DfsH7SROLKpySUbCnElHpeFJbezndiAE1TCicXz97X6WgGjoH
XDv5ogKcQfzScUprVjFXH4jNWoo6U4aVlEgZi5TON1rNwYSR0UqNAOwPVOsbUZUVujncLIwtgjWl
YqqNuFIe/45WYQTriHMOeOXO4Zu349XGEGqdP5tCHZQMcZMeGS/PbCOKEKm9Xj1MDhS61YI3psg7
rtXcvhupU+/3JehMguRZefSI5LKsJ4MziPlMxEsP/ZEIBXablP2VP2HCZGrkAd+3zhRboZdO9bPJ
c42Uz49GiAU15tyDxBceHKbF9+G4fBxGnO2C9g5r5/Mc740UKK6QPt7LH9zZOB+38QPCFpcghqRg
+3bwduZ7PkT9kglxgfxYchExxfomEaQBIW3VpygHzK+qzEqreHL/zv2iAlFXcUmlSA4M39s+nNld
M7bc4c+VRn6qJZLse6dL9U+cpyv21vYv4oxBE8lIzNevlLB9jCHu2XVY1NLh/meR02U+gRXgqfhg
cA8v/dqbODoxI5+s0V7JEPyKlCDiREI241cHjI1Z9C25F2uDcOtPlx5EOqRL48nUMZioZ4ArkTPz
HQ+cbBeDPXQAhcsP8ZfELAiEtAARz018gfU0w9aqOtaunwEDKZeX3wejy9tH9+FytOsQBAgKha57
CS8A1N1jh4jH4bUKb6y8GRWkl/jjx/iIpN2eGjVBJlrVxoEJYL32QLVa21X9+UfGTA/dksu0SG3E
TqRh+trNdhs58TG2+mO8FlJOJiaYgJpuJ7lhrK4+QcUaAnbRNRUVxDjvepHWJQchRR8YX3Mi1OXy
EX839rCDWMewVqJ+VewUfHYQKYKpb19MXHDN/VZ6/6MqZgTYE22c+fXcbY6E+JlodLrbu2fcviPD
WJ8Iqh2+zzbcgPo2VsQLUwfL71Qy59pTRfKFFpvLiPLCmnLfoLfXIMsCdAwms1/WCsoyyidoO5s+
Q4s2jvwmfNgnDmaaUNza/KBWO9pyRE5XV3EmtuF+Od5Cpk50S8obrsa6c6HoMSpcVXEgmu56JhnP
2pV/t21Rib7a1W+VLpEKeGX4a4pJQJSQDkic3gAvLofier1oGzpaTNwRg7AuTAwCBL+ROMsR5UoQ
RKXRXwFuV7H+lbgG/P8o4j+l/Py2pHda6PovgswhEsJGOWd1zwQazLnfZuxJq8OQl5VuFFH39MEC
+od7euMeMjb9fyWn+Nv/hmRaXWgzaHZpXbc4PUlKEjWf3At2EcKCe6umzOLf7kc+bUWz0wifvCuH
rCNbmzrb3GgFTQGBORXs9fRrDV3kjnZynbk6eymnULXi9s+SlFMu8J72W68LolSJw1T5zU6fWxUZ
eC6OzWY2tUDPCFe8A8Vi88L5GfRXBVq1q/bKe6vc8LlKAV67znIXji5SOfHHTvhkiwl/z42Kg6FT
jKpu8SaxiX4swlcyatp917MUslXoIDvEgZEJQcnD+6+dXnRuXR7579hAht3xbKAeWGDFTM0k9mxy
eLfPWi2Bhvhgm7M0tyT2WCTxjrts/RhpZ8D6Si8vjO3Y/w4HZImT8dGmB+Rc65tEI0qku/OpFGAQ
X7JuKQ59DVAl3tLwIHTXueYuDa/mEraXeVqsbva8DA3HkL/OatFj8o3intlI4rGnSSXypj4YrKmI
UmfD+LmXKvolZWgWVDa0XvziDjtrd9fRg5Std2Iw57QDDRIZTUN1ABYghXXD1pAj1mr9Yx2nhCP2
X2FCTd3HrtBA0IZrGoOQooT1Z0BwTMffcV7CxJSOS869fwQgCEykN/7aI+QMCAhjg6QbKArSdYBz
wTtId2IklMQPwBP/IYEHqojNMs+/gd9Co+ewiMgf3fTkkrzLvRsb9LU+5OatJkq81vuMTgG6Uz70
ab40+U9zgJMlAoW1my2QKBdpxloZuSSWmGeVbm+d4PZWudeb8F1MJvAha6kXbwrFCUxwqwlH9QBI
jOP4OiFvqeunRP+/EWs+IPpG8XTn6VCVO3a96cugThHstPatw26HkQ5PRIki0cHldrE0AyQYSwsl
by8YafByjUe8s6b2Nd8pK1hHpF5A3GhVdA42mU4sHHeAsg9Rd0DItbpkT/a9Je8P33/6m5Sb/R6p
Qg9LuPUp2ScdNhpCuztx6t/vrQXJkOsOH8qPLpyeyY1PJaqbh5xppytK/vacofkuG5QAv6Gn6cqG
NQ6ZgwfAkHvZ8d1p/W524LAUO0S/FgXcQELk2LQ/KB9ViI72NOhgHLFkZgNssup0VC0g5IMc3IXE
8SKhPrr0I2SlbzbDZWK6MQnAETofyg9gPd47BySpe3HmqHsy320GSrPSxih1w2/zmIgsJHcV6muu
M9Tqs6oorkSo7U0rM7X44kX1dL6XJb4b8yj3hJTkM6tFADYTAE3duWh5JtxuuPnJ3LnQALJlBkjP
iw7RqWlXa3KHzOPkqsGEHY6MchHwHLbQE+SXwix0LrsCRhqDPo2w+Asm600k4AGcU/HGLrxOwUWW
gb+OR9LXqWGpPgduNfIi8iiYNVXeoVwqwjHnw1by1k0YHosEkqKtP9liRDKJwx7p+nrgy1giprC+
p20W/HT1Pf/NUHm/85FweUdsBkhO72uubGdmt9P+COYyGJJCh7qgh2aCOZVsXCpC0uWran8veY1S
+QDbKFOJ7AcwaXsuZBLHeUZYsa5K8JgOvBHvpI82OpRt0JDFMO7onFzi2fuChEdBRcGcyE6351Dx
WC0INjWkshasmuDhWBXvdRdBFlRyT1XFJs4ZClUkJa6f2keBNJC5rb7vykLQX+z3Y2O9pGMGly5k
SCTHeOSjBDMvZa+WnYJzLJpo3kBTQF/zve/5nJRXFwof/dRvXBM0T39KCARZDJm2oEE3wKBkbi4p
FHcn8xSdiESzSW4XkV2ebIBFc6vAjpInV+U1e9QAO42VusM3QVO5Pt3bhdlaaqx/mHuLbkr1oaGm
fhHJLJ/ja0D0gbkJdAxFeMwYA+KHyvWJW69av2cAOJ1A3y7sS7C4H2+hhZH6M7PnGbvTR2Ht5Eq8
Ktr5/dxViqUtDg4yoD0DrDNgWDfPz+YDlUkz4+VWd1JyOG69OzuzPXI6dibIaraRjVVXpLJ26n4h
3Tn0/lK//pDHpGc5ked5KjLOdswiQsflBQ0HDsXpRKBFRpUiQOTjdRgvnajb4ymohwSC8nZGS4MZ
dIZ0IhLV52ZDuUN/nwpfyE2F7IqMTdoKtA1/vKf/rP1UZdVrCiqyqI7eXg0+ONvSaANQoMNRpoRK
hSkJYPcvjkntHrwq/Hrd9dE80ahUhMqg4Nszx2+AgOT//ZPPMb5gLmeY0NQUOcmMc9RzHr+9iUPV
ySws0YT9d/621yO9W6tUvKW/KxN/TBMAjd0OOKv7f6Vm/PLVtGsg8EvPANDYCmD1UIFQjk0cLC9A
2OaQAHLm6MPRu70xe+1fciDxgglYyMfMMX0StZfYTXNsFkQcT2eQJxxhf+fgjqLM6agAttkWf2r1
d44r8BuY5uAIEF3Hu3scZASgDrjvUmp7phKke6oK2fdsSxYosYZcXAwpjQ9X1szQMPYnyFPg67Ju
pr5VHg/ZoUacfVN13l0gEg/2qxU3uANyxtLhsEO7/ohyZQuu+jiygdchcUl5ss8usnY+MRZn3TlP
TjPCIOxHR7G9hFrvg+p87T8Uv/ilms1qUL4CF11EBfxhM5XyG0Vtj6B8kCdiJolN8BHTucTsllHT
/qPx/G28M/Chqv0LmeK9l1yxjEbA7U9MYig23jc93B3BalVYHAUnjA90baVJxwC63rdKYCti3KIg
Dj+jq9k2MqS4hAr7dwFFL46+EpVntZZ4CfkCnh+tHgkkL7IaoWp3E1dHPlj/RfQGOoXXSw5kdU/x
XtPf9sPLeEGuEDXslb8mpVsC6h66wo1E/1UEudR1591ViN6lx5bpvY3VbWc5fE1KG0a5eedmoxdN
rAPkAuLrTnpkx5mwx22uQ4igbCe6aEWc2TmMBdl9Ol992fU5pbKEdOY5iZPACguttdq/ij2Ag7oF
6LZlZESmIiG0JhmmpJeAsJRBXRJeQ7Qrgv/HdsB3YmDfDIu9FB239zlNQrdrF8s4j2ZIgXBNiEcY
7uzszKjOXuqGjMKLDPaHltaBsJd2y64+TrLp4fV3eWvt45YcBklt/zwvkiQOYo1W2xcLQljXUEQz
rE04FXQM/LkHXGlYoRXdh4fUXGe6sk0p+Gf++fC/eriFjAxPSWdHG5dx3eafRDZaeTw08t4VuiaK
gRPhB8RLtLCh+0IN52f/VvrIwgiPGIvAYKygABCrM0NzBwok7yPViCPMWw9ICsWFqELh88LTf9ow
/gUlKqcv9GYQ5uyigHJLvh5IaZ8twuiLTnjBqWnWpvMwAenwlATthAR/apK4uX/APdhoReztabSI
fK2bimJ8uPKZIpxYNc0hVlU6Vww3eHYewGAngf55hnbsCEygCSlLwvqRDGE2WotajI/9hsqgkATe
kTxU9Y39ElNRmgTg9491POUroK6wL3vszeq4WrkxFCCNyaIoOr/t9RR6piQjWZ4gXL9fL4EPQxRs
qNQ98NwAlBuONaAcz0wLTM6oysWPU7ObzxqUrRPwbcYiopPO0lgeqnYjEYKqT1IzTqvJPu9XKkPU
hVL4lcdTKSK6x7EEEQmdpB1dGqBbj6pb1kk+5cYjciGIYTN8m1RZSU0sVHxTggKQXK3d6qGcaO1j
dVASnvKbnOmGIKdZSpp/ClhUqGOgcJXaa4ez3TqjMzQBdh2ts8Fe/vhze098AVpd2wrGpY8+cdJ9
u1kk3WWlDpelT3denS+FRzHSAHzgC4AUFS9ZAj4jDEclvAJA2U2dmtWlLPsKxzUDH7091X/zdnkL
STIYKrMv1ErrA1MnYbPBrr6gCr2RkcySkYK8ziNg80ldFirgGkt8Cf0Y4XOXWryM9IovUSsKnINl
TV7Xlr/sC1fo20tii2Fd3QCuLTxwd5Dyc3Wbu6ObT/vzp+7zlEWbymEKrvft1JzOXtDjKl/jpNkT
Hm+q/7tBCxt16+Vt6pYiULZJEnlzQzRnLGp0dtfpNNSrx1qjNHFvG0w0qHqXa3vH5hKBrB7kcGDR
uZpAd8IcoBJ4MWKAjBgPZdBEVon4p3qk+4PLy+ygnQchO1R+ofBjVj58zsNWrfKwAJ6HIiS3GKZy
J0Al7huG9GmuAt8qoClWeAKkeO3dlrAzLsYzP+DtDgE7m+feccGd/E/R4/F2GnG4Gh1bz8/YShoS
HHcXIdTbIYZC53VR/iEVJiBdugl+oU+6+IHdCBFOx2u3WAenJ1+VeBa7PJMkEaq9GxhHlyEz4yk0
y5w7txRSxaoDBEb/uCNQAx0W61EISHRZN4V/vEUkuZ7sjPGO6fx1UGwabP03P3/LODOX+4rrHhCd
FpGtkbWn2NEDZBlcgGb/Pu9CUyZk72u76yAA75pYWSTayVhmAeC/XCSDT40hetF3md67AZC4FnWq
MjUfEW0Xi3Dlj4NuCCVlZeG+wk1Ej+N2SKzIYhQ2Ysn40OwKdJS+j9iV+bU6EwxcBYsNCR7bVtks
ZwwRPi+rRJuk/8uVO2uu/9NPOj/73POJBQu/CGcfnsXPYUCSEzxb5dlSJNTfL//dtNRfhc64Aq5J
DK6JKNLV33saeN8AT4XqWZVPRd9h7ZkCjz22lr67ZdPrJg6fTo5Ioarmns+8pKCvS2ghAjtCo55b
6EJTqQY47jnlCXtHdBog+I7xauKCNc2ap2S50/xMHT1E1ToKGlLYbo2Pv+7cK4R1836xOI2o5Uor
rSByFkhAoGfrqsaucXGccXM5qQHbStATneYs3PwVtHvDNWUW5hjN4JF1ySjc4JLm4oZAbcf+bJjw
MNhgMXf6JNJ6OOuTA/22ap4oKE4FVnRA1Ezr8aJiqF0t5NXsSatdh1sjm/baJ5PgeW6W5HpsK8mJ
bWF8oO8A2Q4cwAT1eRiHpV4ZbHNKBeXxUEkO4Q/IlbCvecektK0KMDLp8icrcxR/7lqJHilEP18v
HxaVo4evuHXNcXtHhniw67D4v5Rp5/cP/9IoSGtPp4gWgdbowqVF56LgZE0khDjzK9O7639BDYau
5I50u5A0TD9aON7VUpRiMzCnr3ptikZp1YoWl9Ln5bETNSkfzdvTxmAB/K1dUXvCBl4K7tJBh7/m
0rwRnitJJQv0RzeYx6O0XhMBESl9TvtvaxxE9B7aYDwpSFbCdGqphW8TiJBnt1sCwhaJ9jCmmOZd
CCkm23YB+ODQJLraOjLuwgd7VWRxuJcTG6ryY9P9R6924PWey7rkSztUUC8hI4DF9/bTsQoFVwya
NFQZ1KuAGwjH3SFmM5GqS7cs2Trqg0vK8OaF0FbK3eRdaQllEGF+s8XyKZATTR/TMcxrMTGApCSy
Z/sJD5xAmImTu0TOLz2C3hkJAfM0qzz/e6RcNm5S9xBvqM5Q34D4JWuIO9vuqAh1FLRCSNMCgGAa
2qRCkK5dt55bSMOP0K8IRU4PUf+AY2Qv7xrGtxJkyOTfUopgnwu6I6/yDj2O4jG9DDl06lHbiruS
gBhZzEJhHDP7QoviXai4I+esoYHJg65DUR64sDq43z8hQi2GfJM0/F8+h4YV8DWMKd4kjQsFxHHV
2AOO+Fj8b5Lx/caS49Po/JDtSVTptl2hIXlE7pWfiJkllgV7+f6IQBYvumXhvEKtH20iScZEg0GV
MTJoIYNOil7rB/Bd0j1XEFAo2FhrbLv7OdTwx1XKlVDjvAiFd786/HmdTdlNMqh2EV5GHVc7rx2W
HbUYfArGQfFeA3zFaRFWqFTTBYIbi5LvOiQlRYWRG3dYLeDDdydfMcFD298c69TCTaEVaoNVG18D
RaSB8NIQqvhwnAu72jljNIPfJF0hfj/0ZcdoEf+PB7LEzJN5IskfLaPKlIOknP+D23I7IyPkE7An
sKNBAKh6qASTm56Ugas5GmpRzScv/hRQhpGTxUDBqOM/GFjzj7+CnFMgYDDui+7LCc1B5yNLUJa/
kj+QcwynjNNqIoq/093P8RfbGDnjEwZ52TmMO6Jhm0MLhGJVJ1hX1Ust3YTrrSeDR5TFCxOtlXUL
9ExPUnMUd/5VQxjsrUYhbnsWVze4bIdtvwTXCTdn8q55YQ8/ylMQ7qBld1Pm13Dn2uv/AuM4H1rR
jL7QYdQXPo+cFqJDQn6zuBzcz8X1VolGfL93sX5BxcEXNx1GMCJTAokOya0D/yo+dBcAlXZT1oXG
dHxYWRdC1dj2YtGwL74Oey6SBQVTErZdDi0Hrxfq9DqW4w5nRe0jQbnentxu3jUwfrEJTakLYPLa
qJ585G810aVU8/0Kml4PrSLqbk7ufxVONT7tDmUy5RlSsBRlhSCEl7dEEaa+FHtc355R4No6hUWQ
oOYsj51WdKiw8e7JYQiUjuFDpcemYxiFrvSjz6aoe6YSMLQ0W1hXlPAn9kLvOTNaNuQ5m2RqWJ3G
PobZx6W3hc5AX5y/Qax97DrIeF7PiwuGfsr+oiRAP4iXDRv4i9qJ39q1GhNXYo6YibHOShthZPZg
b+Ao3RHWM5rxR9pG4HKDRlN7MneQMKb38tlszzoPs+yvwrnUG9Ey52OaQO9qqY3TN3Pri8WRa28Q
QtS8okQWOOxayvxUnYRxRPNTcjS/Gn0youMvaJGM2ve1UnndTZpA9dFi/+nqujySEvqiRcLIxAt9
j7IEYFnFgmtvhYLYCT6oc4DTJSUhPjA9w1Z9NznLY7/wBpt4OojT4aWkguPzyQt1zeS9OLIUMfRm
sVjZHIffjMMyNVD2KNv7OgGpqCsFmZuLiE/wotWAqZzMAJoVnodPKAXJQUNRlN5sh0a69cHTOJDT
uBQW2/pB83reGRwvK2ft0NVIz+1yL6CFHZqf3Tw9ykim4JLZ21sRHRP+ik/qq2DWiPUAEci/fqOf
ECgR4XL/prAfyVm+0yMQLCYGhKI+LgITOJ3ixFVFZJcvw312U/1s8kveVI0liBmoHwwMpvLUzx/T
aZFKpa5xsTZ0x68oucF5SUpklDNPkcQ1LFvbo1lzb2fdL7y0Rcj5FGYC2UJOLglMWUzy+7ofkzhR
7uMnKpovM8fdEQznm6BgI14H2VBzWus8Ug1WGn/HyIvHGLhafpWIyEDazDyLd6eakDioSkm8BTxr
KMvyxFZ8cNS6VsDyVMP+5ozgy/9FTg3FvhFBRJsyH5J+tAnftP6P9zESliSZKAW9aTYoEsIRg1om
IhJw3ieM1XCpsF2LVVqYkaI7yneRZ8FzoGqmXhnpmt9sp5tBGQFQGoptHHJIuRwL94c28uZls4Nx
qmrN+U+fnJYnu+xeiYe1RahY0Hws9XQhvgS/W2TK11dB+aP4D7sm3Y4Txvqa5lYO2/lCgsT792LR
FaXeBq74Nb5zU8FkkVXw1V+VcAinned1loIA++tqnE1PiyerxTUjpUTCoOcxyhYZBJuRf2dWHfNh
rgbDzMez2WHkt2kcQzTsAlnWMnzwBizgN4bA8rPP1m0fy162UuzFi19E0ukemzMMXBYBsW1Q/RFc
oBfGbTd3xhaBDgLS1fyrVdSAqyBY+CAxQ0aNfZAqjQBMKIMUtoUkJ54WFtgwJGA3y22VJ5xZGAet
j5GUqbBHKz8oic9bt1p5QqK3E1hnwA2LZrBKMu4FaGu8xbQ6uqL5eiUQMBVoZQWzJrmxlIkmph/e
P5/Xh7tUOPjK5EnuXyceqQT5uEka7FefYhufvWGG3SNQgApewy5TZ0JY8AkKeo1wusRQe/WtgkXj
Ox80TopLlL79KZ2ErtaNTvYsVu9A6Ody2PRjGpqvcRUKuDFhsHKbxQtVBtDo8BAJzPDv133pbksi
2p2G2aDIRBycDKUx+oDqG4eY767kpWmz2L4GInF5zPRQQpV8Bba24fDaKPOsy7yiHNjvK5d+8BfY
px1gBcbEGuM0tpJCeMjHHJPujQMCTb4UZYuzaQONkyIe0pFP+tuuoAkyZo6GO4A+0V4FDlkyJkF0
oGsCh4iBKxXiCNiw68VSu9ozx91z5hszASfTxBm8Q9LP5FlsRuqFw3fWyKxF1UkH1ub2WhuftATu
R6jz8FFyIs+b+5++2NTWUG1mcYa7hjlo60YL9dWHBTvqy2EKUqLgPLysu0FrPg1jgfLoYAT/jADt
LW1T5NZC1xVwLXjmoltHfZu+3DY48EfB8XWBepLiuPki9jzxpm92/HHL7H9QB2dLNDP2FkztsvwI
nbttD/W+EbuSCIj7ytTVH0tlX2/0O7lqhkDT9ubckDiAcamAxrzZvThlAy4x4KX4RvmkOWkFy17a
JMnFesCjvkht9C9PupZgCUztJG0j4pMbf4DByiDiN3Wg9cxFohlocTLi9WyJ3jIiW0EtsCgcqLvN
9WuPtVPjgQ9IEsIlFPlT9uhJKFwUukgEjs7T+CGud3UNLgIovFka9wrOpQkVtVfr39Qeag0D3DIp
oY77cLoPAIJwiPndDcXwu6O70zY62XtSqhzZ0cxXE8I6UtZiyREUV3vR/lNM5EiWG9J1wZapEoag
g34uOu/gD3YifW81vWRj/Kp8PoOqWUAFC9J31m252HWyf5HXDd118yc7xwYXxrGdIVWqtPyXjiVW
tYfN+5JDJHkzpR4L7WXDXBYRpHCvgacAQknh7dLmXc4cUcal4OcQBLnKfLMLMyGjGFcUios0RCp5
UZrpNICLlk+vOYFS/9hajMvMbxQYByTZmcZKYBmN33i/084Q2ZdMWzunQVbWB5RGA0FD0bJk9epw
tzM800diS8Vndhkb+4JQhnnYkvq9tPDWd/Yqot1XvliUE63m1x7Pg/YhaH6N2iljP3fSWOIHMU/C
pFOO+EXZA1rE8mewN7+cqiqJFQokU26OjzHL5Z4UXtBRMscIGJsOrSWZfOKU+4gvLe+FnsHrz1Nn
MAEOMjBZzMXrs3W6A32DPXJ2pnVFqTZNSJINhn0z212SjErHGq7BQX6EEVCwLUlJ1nOPeWPB8MOG
ff64MZIBI3gQO8uEVotzhV34l6AhijGE2dxK/9lhiFpNRg8TujiT6zRbEWf3UXA3ymVnqjdLR+rJ
TOpov62ceYIofDTv138/Hncblj+OOkO+cL6wLb6CPMwfWsoGAi7EZYOS6YoEeKNNFlCG3wV7BUVZ
Gaw3M0pR8uyCixSVp4YJ8+npyVfic3mkoID7O3oAu3igLW/3vBQiSOALAzHYdvi2x7FX20Kux+wW
DCx5E726q272ZUZ96L+rrHWPVirK2SFQT7Vcoo9irlkMhp48yrGwP/sJb4oE8TcLOVrI8ifhvLNj
BIdinVolKJYltLH3vPhhmul2PZQ65Hz95aXZ25exAaW6cepMcVGHeI5ltYhnwCYjH1zpJjyC+AHw
8cmfC8+Rc4lO/wH9+xCXQmvMZ35QLhtpMjeebd6OYUDo9zIxaofM6LIZrnpmhI9SfyV15s8fmUfd
/VUAbPOs+c5/vko74gBEDS7PEOcOYwbt7rJy0APeO7tnHf3P5tHEE7TzHDwl1GR/S3q9SMYoNvkz
umGdTc4UfwL7GsMIKnOncu0QC+wYvr321kopPtSrc+Ln9FXHhWXzQbJu1oixsbqCNUJ0qMimadCu
mt6icUvvA5WDzRZYoDyvV3MkDyNFuB2II5yP/HwKoLwivjC0hcUQvkqQjyQBJGP+J8FlWIreiL7d
9q6ch5xB1d6/I7r31lh2Xl1tr2c8LV62WZloW5eAq48KzVH5R8pkAk5FoWm/6AbRdwpVt6L47/0Q
hq5G2ICw1qbThHCwcripO0R5iFvSYdqR0Oen0Qj+SVZp1l+EvQ1Ji9EdnM5z8IrFt1rPFb13LjbZ
ubbZ9rq/G6PsJEhKrSZJgKLWN86CPVBq0+iGwD4Vg/KmnS+gVABG/dl19R6zcO83vbvLAYLaw8AR
SyELXshcKcDrO5q34CDCzqKySMs6SvawCkYWMw1mtiShSbDEYutZSTpl9ztE6gfTQXd9BqYro7kx
grMeNT1e+NcNREFqm1Hbmb745/HIJT+scs6bCgXbSB14dNQ3r422hEVHB4X4zGTprwpgb2rh4rsx
eH+zE4+nLukBh4ws4NFmPb4tfAwxm8F21G5mgtoBp0+g1vz9+k3vbtKjBI7uNnL35NmxgES4FSJd
xZ+NvDMq0PrkLFahK970r9Jc3CqQQ63d+xp0FEY75dx/DxEmdNtZNWRa1yfMp6ZCPc3tTtFH0qmo
shyYeJe+iD8Zqw09oe5dDgTe0+b02QWIyEs3oAbqQYS8PKcHX/rvN6RaUPL9gsMHdj4NS1whrXxH
ASBa6mHLBN/WlbCEFm4LGzuW4wnSV8Z6JhMBzLm0WNMTxhnemeRTM2z0VR/2gjLlDvOjIENrK5Zg
BPV8835Mgb4pNooHHWVdLpclBKxB2USf+Wo4tE/6YPDh7SteoV6MUjgML7BC+dbLRi5gE7008uc0
jd0CfZsQY8iO5xB53GOWX+DHWpTpKraLAKK4MFfqzyi8mJa8v+TPzEs7FEBJ5ZKuofzVGERCQ6oz
AJj/ePueHjp1htrJk8fVa0sMJO75UUcuM9vqf3gBNxNGSWhyofYc4aER9VXrHcZBukyWtlEIB4+I
YD5oP5JQz6vBGmwmmt9AceXVBEJk23GIiSggKcjl+Ua+QU+dc1osBK0QVhdNTax/R6DhKwGabzNg
Y7hJ7Vcs9Qa9JcxrTioElhMMIPSpm7YGqTU4EPnvGXyGaqFsom4KBKJ60lPK7vjzYwQx9y/2poYi
c50nPivRv5tO07xw+udGzOHiySxcmfVKZSe1jCa80R4agnmyC2ZwsSGMeHLynbTl6Yfdg78p0qbx
P+AaAiHbXACXWjqN6w9b/lPl+sdLs6DGm8T46Sne3dV22PeW72QYtukh26LQfCO2iPxgURabiARQ
LTiTiPerWtAEuYXSw1Nt9neMMuIp10jNpZ35+MXHCva6R1ypKfY9MmcSjLflfAkL/Y5q6vj/Jmc7
m3sLroJQ3IE/eEoN2jgKB+bszVoDFkR9j9lizZ/k5rOtHmcCSFvnsGGCUrDPPI/TbE4NMpK+4Fl5
JJosLrY3nQkLjYYnX+bb+BABzVJxxa9LuWrHSatfy7mJVRqEHSg9FYW+PLruQz15fkeLoQzuyfAn
/EZ4hVwJkYXPybr0Aya02c9brg/OE6W+fRfBgzH6hJj2fzy0GHttwhwYzpwm5WEBZF9p2O1vRKyr
akNiGhUeewfg195gfLM14tyM3s2yb5DYhNPo5VTj0eqTkexE2xw0w8hachg7J/QxGv8o+cHhbSPB
zTe5+9Nuf1BLTRilh0/EymnBc4pF670V+BLGqp2p4CAia4ggeijgavwtRsbrdl8QGp4liGG7KNlz
5WrZdogs5PHFscZgTooEcePvTlMu8ZjyqC8oCLh6mXXYav4h2WbXwtXNjcVUkN+zmKLonBW53wHf
RIDHlHlToHxZk1rPBUSuB9G9HA5hHArq+bldg0iLFE2LPRiMTSo+N+CXXePnxKS/yzXCb6GwQloR
P9t5PZsixP+iGxkxRrbFrgoXOcCubfq/bpVV/8qbMLmY9hjs5CFQQXQD4ReNJPOM/BRnfq1PeGLm
ACOAAwD4+xlSjtfGqR1F6Tc9usLaVnF9k2AY7/+Qdv16rEeKxUKjjWVKVAs340IQWk+fW5PUQoi5
tbMMJKIQ4r3sum12z7GFIExWsw5WF/VRAvHn2zVywnRLVhG+tz99okj0+CoF6HZlU9yvOMQmNpRr
1aG8aRTzNC8gpYACFxxVOuaLs1+bxRnFKlko6/ZhPkfWI50XXI3eDTdCNhaSGVQBQPy0TtDELkw4
oEuUBn0Rm/w8PIQYZt8yL4/6Ex3sP0a+ouNnwtaJbvY29rNu8nDAeZxw4uNY3DKYC3FEcsTKbBP3
fLqSYru8CCqOC+x+/HoKhXVRZKiyXep2AqXnF9KqeGlgwtISlXd/JxZL23ZNaxYxhm5woMGh2bYa
TEDK289SGqq36hgRAL0t9Pc7b0XXCinq2KGLdobMIuAL9gSwzC8SPa5XuiMhvi3qqrd/zAZfcM5F
RdEZTbBWN1NJA2025l6IhrYBSgdSsAsk2tTX0+8W7Jo3xvUI4dSDoAXGGNv9STLkJ8skQKcAYm91
cIF+TnXHji6GZD6nBC0YwOH6PN8eIYzWELcG8FScul+MZvCctGZ+jZRk4FFsuf4X/LPD9YtbaV+5
dQ0cQ9xfJb8YTY1hTWaUOx1mInTaA9TZ+lmcCrgLvqqZ+nAcXr9w4g0tKGfKYDBWYnt+geg99x4u
v/SMJ1Tmjfeo4YhP7H2GjDalBvGMUzzAN0J0F3CM4kMcfc+J8mdaHsl43O6vrhuXMTa9omPmsW/y
Fp+3roK78wLvF3RMB58W9jyTvfoCUKJ3if6J/gf/UE7eNZIpGcg+uTEGkCvZLwjhjTW7faO7kz4g
oeguVf13G9f+U4xvDVU3vfsnPK/wExjQgylIjahcNVwwhOb1Bf+sFpWAXeljVxVIlSHO5c+X9V/Z
MXrE0Pssnuj2JDOIJSXewekMBaCwWFhrVcj2DKUEKC/qXeFPlTaFIhbN14ilUdnRj17ZZaeHaJVa
EwQ9R2vjo2grcKBRaQ1dNlBQEHV+7iwXj/HN3wtbqbynxO3h9eiIhKnVi4ZQT7n+3D/s1VJfJ2mB
0GvXZwPL3oIJ2g5FE3Q/Xeh/A2zVyiiUYPn5IVPE3tBZNdLXGHFmZUrzCZane6tdn+s23zk9dnRQ
k6Ie2HjfSU0/soXyxhA5xoc1lbXwzdRsrQmngN5oZ1I5wtLoe7KEMVF9kjTvyHM+pvv3XWZp0J99
LZXEjejy2DwH62vnCs4+5FEVZp5DUCyYA6kBhVQAWwaOlJTGGw45VqOiuJvhCEiSBSEzoXLGpro7
5VVFBXnGhFImXlieGQzzkG6frItEhrKw8IhguaXXg51hes9ocabV+W/QnTdSAKp7AsXohO+iBEKl
6kyGHQz14PI5V50uB4GD36e3ySkITDlZY7wtlAMx60np14fmG7doenpb4wajACwhjudzqDXXH2b9
9XFcz2zIEUppmDGOMzIVWaRHdyrjeIx2VYURcCiYNhDkeYem+IVXN6gMtlZWC3qxXG/OhhYknBQ0
9n907Tz6LBxuEL5vBbBlJAAcIre86BxJfEnDcVHtVBKtPD+o0MEKtPyb7ShIxzSxqkJ+ZD/GebPo
O/6krueNef5h3Iwp/bDv1sh0tqIx6IGBjQZSzCeXhFTdaiFR0nNO5dXHG+L7EAX2spsV78uW5WnF
Z58D2aSCX0U8JJR/olMSf62GAe5TRrdt/HeWgoqVvJBGZE3Tv1HvpigVF2Hdxm5TyYMwOsdyERSl
cCpK1ZDqfKjjePY+Ilrq9DVXwGzQh9D9HcHuDVzQKnBEJRhefrHEm7WzI/dLuxLAnWbfObtfVOWe
qY63f/qCICJxqOQcWe9FY1rVqrmqMLZHygVf6llA0FKn3iiniDUsp7cULR/w8LIqQ8T/JKKjAujR
mGZsbI1Ua2eU2tONwQ4pYQFHwOdF19VIxwdsj/TV+dRbuCp9amLWbSq+J627/n89yKyY5pu+ZmD5
fWCtFtkumtl5S17VZGAsreV7JH5kLyt3drufektR5Mna5eCzIidyApGK4hQ3oMwiH1X55nk3GMcX
DF8DP/NEXJhfGWrG+Hd83oV+gvm6fQKQjglpWX+qGDFUey8LCGfx2LwAtTj65EIm79Vk9AD6+VzU
psqjSjSLOpzDJTXARqj/NioAHcgw1GBw1X9oDRa4gCRZPTrqkPHtNVTYzN3jYt2JdknmbPW3uV3s
qihhlIimG+i1YxahB4XLMQtVTZ1ZLxBBmbZ76tMBDN5FbZsPHW6P+ZL/u8IZpcrs0ZzPEIX1n9v5
YEZJnurc2eUUsipvRB1sXcgSd7leBD0+/uj3qAPy/nBNWB4HrfxlQotAYO7GpZm+mXXFI/GL+Km8
XsRHaDaauL+U2h2l7zH8SRIUAGiWtFqy5Q1riQilOt4XzsYWrsZpC7rYH9emEkZLMN4CwsOV4vj2
mSRD2lbWyWIfCsILDqAFUbQpW+8J6LL85jHGKMk4Eyf3JOkzyoGabj4ta95xjIP4f47+ReCYJLTZ
I+6WOSjgE7nRKm/VS+gj5QcGEd1WEr5R0I9p+M4SS6e3g7OnfP8gRrYnALcZPFfmnVXVkw0TIJUz
Bizkrm2ZodTwNbK4i1jJy6rQW3CUhemqQtWUyq0asCjhP8o6zIpN0wncmzZlhUWphLjwcRQ+gzag
yzFkhK/DHEVgk6MSoPrNkx1j42kp8Hq/dLVL9wAfZ77Z63tG7sDEkmhrcMh0ond4qvYOl4JPiMBK
f106S5PD4WK+ptbV/aDrxSXMB5VX8TxTMj+CcYAy0+fq7pG5yWWPSEcZI2D+g9BWqtKMQCyc3W3m
Fd4O5T4mJOS/p1ccj3tEaiJWq6LaQpdeKB3MDEqxeAU9K17dy0Df9ZSlyrOlVJaDIp62UDnAbZ7y
tJvfz9L9L6iRMDTbQVeDQ8G8/O9ArgFUJzU56GXOcvPZPakk2vBGcpc67qn9DQmp8eqfS1TxZhfY
y2DegG657wm1/a8ar/3dQYFjTa8Fm88Qqhx0Bi4jlYVS9odOaWJkDA/ggj8QnoINKd8VN2Iw5/aj
uIpitWQG8fORf5BTmEQj/oT4ZvLltjykiBTzBKHxawsovQj5RlkFWIcl2btDVoUa0EXxGva2aDn/
L4iDyNkehm5ehEcki0dVMizj9+G0+CadBJPmsEuA4BwFVig1aKd8UhngS2YH3Xw0jVndZXjjhGPA
NZSZetlHNAO1DNv48UQmM+N6+IUHEsCU9C6UcB9UbSPPo+2stZYtq4mv7vaFbjLKXxxPQAoYr4tV
crugCnFu2+f8CyROQODGGCaGIsSQi//RlWx1OMybGXpgf4mNYvMvygKAGtoLlCKQlBMtfZ3deMEt
+ztaj4VeqQDx4gs8cwUBrymuVYxOkTqYJK4P4Djsf3dAFrsoD0fUZBvgGE9wLNg6kbdJo/3ZHpai
sGZO3F2sVccZTkY3v21KUvpAD4MTf1L1GGPzyYu+Y5AO5UWO1qERrDkfEo5u6wz/sMDVbbZWNMVz
5QFVkxb4lKIsp0/eXKtRrkDouJZuvfqAMqzFHM3Pcq2kzGrcqgiHUmfUCsY7gAFWZqn4trYtVe3d
a9x+Q7oI5qo8VKHDOfmZjaGZURFMSH+qemEbODzYEiZPJmZQ5lT9ya4GqJhJ5N8kcHcy2FGqdW3H
ztclkvDcVZan/Nn8LysHhDdPbcmL29D3gC2jQZG8mOUW19QwSfBYgG4+L60x1phgHyX0FJt4dGOn
uUcjsaaBtOTtXp4zq79sf+1t3lxlB3hDwUqFhERBAEbAUP2ZTVe46Hgans/H02CuRqG2zb6b1Bk7
SlkqaD+89iEBvvBDXDjUXeih4LchUqipLpbJX9BPk39LwosT0NOxIvthnJIGjAp87geNo+CsJdZu
oqfkjcV+V5HVLqpS60zhru94QEkLli3tIcUvTQrVKxNhr7LD+YxrPe2rnJnt0RxKwjaXg550Or+B
x0gJy32BmWgleR5+awOxZbxuQWSDLJCpn5m8huBLcO1pklhuXfYoXtZBwB7aQCotaUwGhdlvN7Bc
mBNyBe98vmAa3jOtL3g+AcXo4J5ViqOLymVzvHwlOLn0w6jQbxaVM9zh4Z7gP5pMnp4W1uiG861U
UC+9hbpBg+gU6x7/cN4VQlsYqmQsl1+pvsP7WJAZcDCTlOTg7VqNWsoErkU3qOalAfp+d4nbMO/e
M0JCQDQOZiLICKN6b/Lar52qY9CSs+4TvlxUpDHzXnCCcSu1eFb42n/G0s6q3ai5KE6tbFa1ILF8
I6C7EQmlhcEcQrqPDzip6ppr5Vc49B+GNAjrF+ePTCzuuF5N8YWD8JxfOHUTJfQ17zeOfj1VjON1
6MmEVzKPldac0GsnCPg6tgYJC7287z+OJ2iHuE7bHZt9dR+x6J2LAn3eT3DOOIfdlCoYefhzX9Px
ANwpuRNJmRjYY+kMBO9mXVIso3fNfYFh/QRANDnsGtGA/s1pnQeRHHmNR8jboEcG+QWvEKco7BzM
Iv1DQ7Uf7V/1MyuSkW4JskH5cHWxcCmfk/XEyjehoaKuT0zF8sRhBKvOvXrFrBu56n5yTHjGd7d5
lW1VAJyA+4g7gaNKc/t3+jNox5moEUMOF63lF5Qiv8EmEKNbb7GiQi07dz7j5OdMBxPfQ9syMp1v
ekCsBWOe2JA8e1Zzh5tsnhIs6tbS2UZXtpOGZjKPXrUwqwRj+Ie1FfJoOccKlc/n4BRCJUECaP7X
pv5G1BSgIROEZ5KjkmAhsnr8mXnr/di2mPGMltg/AWx0qvgoxIgFrf0xEEDYXsKwF064FVTiZWOl
iScGLcv7FIo5qb1yVYoA3FiV1xBZ6Bo0ccaATU0bJFLCvbjzy6TI/xeD1QwZDixGsQ5OXCHPDssB
vpGL+6bM5dMN+cVmhgAxBF8lTFaoz4ZVFT4VkCKwMwiHBm6hfWo+21hfm4Z/SKkzMEAQ1caKkBEj
qLkjgdmtND9ZRSt25o4RLDLqkTiCWWHyZSsaip45txrbqLtS2tPreVbCVUKITE/0htd62rJOUXdn
jWuhBOBp9VhqF7dEKOcxuhC2i2D0SCbNUqY4fBHou81cdr8Nj1t33boJi55vC08bDKIldCooCGj1
toGTnf8GuMi5NVPIp0MlkdtKPf/DGklrBtkgSUGNhvBosDuiDf/DDYD2vpmGsFZ1eagGQ/w6uKaJ
Brmp2BvtxBIvT+YB8/1w88KmaARzklBZNHeRbzHcDfdvvelccTj5Nxk1BbKyUPsia+2KuNrPtrvg
kKc5aeuh3D2XP73GYX3I5j5t8p8LSTH2jpmn+LNmcJ2UDDpGqvxyyRiybWrZnbBpfX9Vjy9zt75D
Jhbist2g4ouUx8MO7VFf2qbU2CQ6bcMkDvEkm08U4+fUz5CkYFHR+ZsukWump99rskc6ZU6dd9y0
VlY6SfF2awK5R0zwT4SyWLnevsD+eej65MHXElj6SawEVizbF9fAEaSHeZVL36BoiN7N8TkPlS1U
0FdVWhB2HR66JNv5ZkyyYzGP8uskWbIIVqdlgNRiAWJQJQfJMpKL1+fRRBqHb4UmB5u//3OiFCTQ
zrBT8AJp99zKy4cdOm/ItIkVQ3qOnQiaN99qu5CcRebx39OUX3VSIAewBWJJI4feb7VfaB5rI05A
3NjHmVOY1zBDDAgqJDNgNFaLzn2j8VyCKkT/0AZbhcFi5IWs37S8KS/nmAe3xo+FRqoz6KpLJrqf
c0lWgFwN1dOJ+XcFw3Vh4ZEXWaHxItFxAaqpY0Ax8j2timKNkAT9g3Z33/gUU91Prm1OTe9eaNyg
LGwopbFX/ZbD26BMZRXEOuW+aHBkMzJ0AagZ7MDFPfvT7UFAZtAu/i11BEajeRb96ejOWrrGfl3Z
Lrd8MvgpslDvFj3u2ct4pKtMN1hldjjVF81tl3SZ0xALWUj3N52fa/gmE0af7Btch6tJd4CKCwMN
+2COhN4/DTZ1nsnWjyeQQi/iOMG2rqPhr2ahCwMOFqqtotffRnPKfaNQhAtqxsCEbIJd3d2wB41C
JGbGrVYgkGgfy72mmRwcG12rVm2KJtyZLL6jEkOI7ES1luG5+XxbqwvblaYPh5zMemD4F1hDiW7C
8CuIMZlbA+ktf8zzF9hzklPXBCe17EI3msG/kvwcG0NkmsTKRcTmn9aUe1Nis2wGzPv0JTTyYAQi
86zXZOkFKSS0T/cfFIceHdzP9nDYAWDDhljJprAlpdQC3LNxmH8MTts2X9mmibu7hXH32X6sm9x4
mfSJMZrxPYkF7MxSnhI7ZYA8iZ/WP+nKi1H77NFlVUByFGDH3x4S5IQZnSAwSgnGNqu7d73eOKUQ
8m81K5Hg7WZ+04upHK4iYn/wwHjkXxywWKLh+GGUXalQilNuIiiRWg53S3lbsgRGy63FtTrZeYz1
rpMMhdIAhEpj+pKyS5UjjidNheExSggY0mWL5TD5x/HftHsLW3FE6gTs0gXxDmZQsRFKrJTsjbc1
Wmpgdk+Tkwfs6ySEURWq+G0Iorpx0JmHlbZBu2bZKTl69ErJm8kOrqHLCkQMrMNTwBP8LKDHfkVA
3/BJuzc2G7DniXSSP1Ej7mVBLIvHOCC4LiI1J/ujA8tj3EyJb7kvZ+f0XXEwYtmblrid487Idhpz
jHDbHx3Yisw8qxIcS6bYhaiV6fFngXqTOZ+BY85K3/t1lyNBzWCLPsmmSwIYYtnrbWRI84dM40sM
gvXfo7ExNUM6gET6ckgi6Cs06f7x7jU9Y9hdF1hccr/aBKiKHvQ7dODdaa5HQQVeFix3QZ/nany9
kX10JMKglu+Obpkhtz7w2w5kGBsYQ58Qwkant6JiafvlY+8T49CCtof3LtIZgmzupHI42RBwd+PZ
mtkG0R7b/Ulj2aVdMAfvhSpp1DsNOLiXSe+BAw4PTIvq+VPhdWNao+DQhOgLM9c7bTtQ0efN2EbZ
j7BjXaapvJkGReoHmYx8v4OT0nfOO1X5x0LIcby3Rr9YcdAagVKbhnoA1woyFXrsT7kjhnT+6N/n
rDQzKM7tdQ28M2bffX1hCxdZqpk3XLfr148UNg3GLcH7axtn4gxdMFiNqZrOOOi/M0Zg5b9QLYhv
X0W+jQIchx1/51ywkb1Ed/tjMc2nd2X265F5ZTPN8qQxh/N8HlCvtX99zK/y2Za6bGAo+CwJ/r5O
zjqEqerljrWT+YGbCXAamnusZVwvEEwgrwHTTiMdDGGMaykN6N/sH/eOS69R67E8iJxPcvLs1aVQ
SJ58e/0gYbFF19DzdHJfedhM4nn0umbY7II2LX2olhE1oSoGgYi5QLiCXAEH0/l+ZgrYrvNOCYJD
TS2VE3y78t16xiI1sfwKYGf1Eolm35ee2dYnbq59ca5qehtel08SVi2JZcmgaxWpJnzrWDpWuR4m
Gs7bbsON89LawlgwzhB/Z4pSPLm93e6vm2Aje4lRRTDNeb2mYFOfSbGwX/2THMdVSUy4Gv+W7N9S
vkjfnZSIpRzrVIsIw8xY9Hk2ZX7nKmg2/334YYVs38kP5dyS4Q3uA381ECbX81K39SvCuWBzwfDd
XrJblBirQ4ajE4rEMzFijRemhHd5xzB/H7pZO4bzaAJYTq/Pz7w3BjB5ZgQtMCMDB90wwa4M1/p1
2+ky6eXH0ATApikgtLemClw3UhJzuEXd7YHU+6e9IksTjYwv7PNQ3AaQYibveCY44WP/AbuBGLwk
p4/LmRbk9CcPj88yg1nHsdlFoDCDD2F2QUWQVlIOU4I/HN8+BOb/TF+JHPVwaZ361N9Ancf21iz8
ye4PmEvKQm+QC/AL1iakuDZUKJG+JIq1ww5lkNxphhP38uOm3nHLX3L7MyG20BfVcqXwx2KFCXf1
r2E51x+PxKQmP6cZwNUtI+5qc+GG+eLzO3CI2uWY0eYPcaiWyjkOzY0N1x1yun7S+fM/ZoPn3SJ3
m0cAPhZ2XsMJTzoj9eMmU7NeYr5ATxy6QI8SNFEAKDIx7bPmYIeQBJ8EHxwdqkZ2zBy2+jFJa+Pe
q0NLn8PiCq0KWBIiA81IdLnU+2LmkCzMkRgH4FNCLI57orkhKOP+ukypaONKdlZmGwDkKSBVfh0l
KFcIfzKqAYAawgbkboYLH94+3vbIuwjMp1zgVuvSpQMYO0YI1HaNPeSZZ9t/zdB4pRql87v+LBjL
vkuw0Q269Rkulu7xx/uttBtuBqlR2qYJE8B8mB4IHFMvzxXJe8ASVIhDwlfZ3xz3J+LpQ8zVH+1D
PTmWCKa5W4PQ9LgyZM9xAaRhrUNqhNjUd0iSorFDSmbXubo0Y+EKu2uLuyUfDvCORPjGcrbLO1wI
JR55lGMh/u0/0Q8Xt5gwNMzqJJhN2i2uowQP/MRPEPzfaWjcXPOSyMAelGtSYobReSQ1wumuDggY
NPH8oYTndQt25FURvSbeGbv5cZuNI1RG57CwIubXTs6Do8d5HVBaPP3tyGwKLbCewrn/X8DVHkDW
2AJ2/IG1Jf9e+atE1YkGhn2K+Qhgtyws78w7sG69C1zLXmrsoXjCK61DxLI5UwsLWm4c5KlV7l+W
zb6w8wz7gOF8aZP5cK8ff88YvNTK8xBZU2n4GEnroAp5kD8lWndPhkTSQwBeqeVm/OUWU1dgo9Ov
QEBCaOINDzEy8fdhAbRN9QIwJ4wPYBWdRYH3jrTt+188sDwcEePnJmeFz97Ypj2l4iWC6Hs6L48i
RgotVtebjVfdKTmCZu6AGRIgdo4V4e3Qx6hDkOJiLgUAwpX8El9kfDlRPd9oMVwqvQeTezzMabCi
kTHtok3ODXqAY8mzIcfHSg7TmCkqrlaTPnRefONtf+1aO8AFuGqfgFR2sMaye80epKm5qYVzx0J8
w5rr5QXY5SIUqVtznrs8UogSY9XYk+9kya9R1UiJfrN3JY5Zd7eUXPOUQ+EqwklViHCVJuEDJMPI
FyFVtoZHBtBhc9/vBlYIpPsyLcWDGCmUxP3uMkVdz0a4pwynjddteew0aXKdfqX+2RI042MQzBJj
5UAMgkwLKQyXjVLhA+rrVF8pLSf7DUAFwn5s0K3+03U8AEPXGxIXsL7dH/YK/09s2lHoctX2Jr1D
Lxxy1uK0oi8kncJHEkd0OVt7JR+6Yv1v2Bj+H9njnpUg9uBfNRvKEFWKp+MNjNapZ5/eo75HRmVJ
XkfKbWu+X4efG0dxoagyoKm9Co6oa5nOm4lzwFhmJ/9IXfpHhA5DzxHz8M+oJLqZ37oN/Koofgg6
PG5zhX9Pz9j9wjOvVOPL/vsEGCyazDubAceuZgq1phgK2SLop3AS7WCMdvv4FS3toX1WapwrriZH
m2H1+fuVhEEkUtFMj6WQE7xW/YfqHHWb71y1VV39aie/AF21NtUWFhFWXskiiBbP9Y/wCp/zchW6
xaNL4SgvYTEurS1tkiLMgRKjygxlM29aXPKCJT+BpgV3x6r6JqNFIMcRYJUIDj8fqaVC2kNeo2kr
79tWR02J/NPbvbURR7pEAHHJTtrUgT8GxzDiWwCHS1fK+suWFcrD8M4Plu1YyLInuuSOVe2/yJLp
H7zjbWOZez35u6uM8EzJFZaW5IRCUaoj4/KozArbXPb94kXTbA5bRqTnCc9wHz/bkT7EW0l6h99C
qSqYz+FENnaW2Z0CzcVq135/h0jtGnxi18/92XXQOQJ3y6i9rUQ6Mq1Gh5Qu9ZZFNprEssTJsGII
4XJ0ewYGTg7vSx18A1fdEJKiJyz71ULrLp+3vZbmWEbsioPZ9PV9A+6outhWscMbTZXfTcWDYzlC
241rKZBeqG+rp8c+MazOOjT6dwG32vozRk6AUey4MBpyuRm16iZncQMRt4pKRixsxd4fm9t1dI7Q
ty3RVidIoTUMKJ38kkwDsRYvithyJjSUU+QS0LE9qi/hWhtf8haOwKnjttKVONEroOF2ZlpyVrkR
13TfAJVB5hM6zALV/VQQv1jQfpgeHmZJhrjabgX7VcUkTDy64QfhAIEdjDmq7fi+1PNlrhpwE1wr
xGRdhJcu/UL+IGJpT38p1VCUdeuR3yp2BoW//uh/xeuxp4amCO9Lolg/ULMl7oNPOWdE9DyXpDUd
Wt46RXFuMlLuGJ9QOxwLGAnfTjvIVRUquFyln8/mjJGaH9aAldh03DflB/7UcYpfmROqtn7AgLEs
rAl0lPatHaTiNdU/YaDV73Pr/beHtftHClz03yxU7n0PmIVdJhOzuBJ3Z7Rgt/2q+SNPERgs7nCP
fiDs/6hdH+MJtq4Sl3hS0PyPgeG9SCi9N0N0oxUbHDSQaNzh7VJBgqg97KfqzxltE1qv/RJ1UhAO
rKyy09Hvo1h0tknpmof47UqIlbzkCCS8a7BfV128brTxWDtSbxnH/CCTXT7jUsS7f5EX/PaMkUsb
EyufewfPlQgst5c8XcnxqdP5DjtXOkRGEEGAwVxA9Z5yYUcvi5Xlbt8gQut2Ugmt8TowV71fJ9Xz
hVfI1G5I1ro9cFOUnj7QxRkpKEffH9meETdKQbwa/kar+0/VjtHoTCseysu49D9LBX5EGg6cCxVi
xIr8Ef7lWSgTbkSqPgXJb08surtozFlF7bUcOts6k/fEsymvd+ph3x2BntKLuyn8cR0NPKV+4zbn
1YbRYTJB8L6HZ2f0VF9+X2Cq80939fHMwJYcj3xoBb8YbuVtODbsMXR/609ZWGMexSu43sRagmcU
a8K6qkPy2MYJfEgsJ37bzb8rEVhOWdJ+0tr9YriIJ6nX6mPQR7teJfgdsKCp2dA+GTm3myiQ9qJx
dGScC6k8pk44aoL7D5Zvkd3NCMS6rpB/uiF4CKkMIgiGlrfN+NkQc/17dVpnBEIE9tr4/39aw7g/
ZQxzJdZkWzY2n1mRHfZNFZaYNP1UNLDMdjhJ86H8OcRETlF93zTikRf2M7firTOrFMo94g+49S08
mGuUwfK8RRZbfRzS+tvIh/xgDheqcGBetUjQMIr5YOEBBn9B881LL841sKmchmJ/zix93XbohilE
bJzyB0ZqLG/LgX7lAasQidbM2uyTWlzCnnWpJ4cIz1mia/+1EjV7z3sWO5v2D7AQJPPULe1f6/BS
IrQqivyinw+pjOAPs+jcwaIRSNC7ta7Eyao+lgqyVyclx/abuln5EkdBompbNt+5dyRMDrVfMx4f
1TFgva333V5xOQOasEQzybNU9w5S4EbWw/YP4g2Le7cIkakVhUE8GTavEQN6PMs9a/NXUx4mg8yL
6mcksm+KQHf1GhQMEZv+JiOpGRPcvrWUbUD+L3DmjmwQtynbNgPZILD02dD71ckBjqpebydcxO0+
0t5GnYhF7sytKXSGgVq1EzDt3d/PjOgUFjzpdPIhFGTTSiaqfBKrsy8wClkcv5SarvvHhaJ8NTwa
wBsmJutaN405cQyywyx9gr6DJ+GdY+FySlX4mEpBKVCrh2iSMVlrUdSiIv90JZVdtg2Uifc2eK2R
WG7gQKlIoxNARFIz8CErxZ0ssLtRl4XsOzmu9rbcZFqcv4tZ8DA0UpP9MetXanTkMeB3J0G3e/H3
WLk6xNGTh7KiSTXv2IYVDcZpZrYtUAZ9a6NCE+YMPYc3O0LSBwp00bT6QvBwlU4sxsyNsXWTM0lm
9x/CNk61GYXbG7mDeHMZ+wOuBwR2jm8EvWakSrQNt65PJ/JO9xU7mIUyOx0sy8ZWTvWLdh2mu/jR
owAB3VDym90t0wXOt0RJtV/6cWwC62OVzUqrlgWdrP7M8+3xGofNk0HeFzWRrVyBEpJITcCkBnNG
wX4LKU+AnPT385qSDgFHbMnCYWsqfEINshoiPienZIW9HJXE8RFlvr8iMIyv96BNmK9TXoTJbDm/
5IttWz2UxRunrK7X/NGqHnAZ0nb7vAjFPapdw7zX7kOPqWVHu8pWOc0J7guQhVXdNokP16H08a3T
WtKLFFUsqmEvutAFwNeq2CPNwmUU698ezcL5Z0IZK0kTtDaUz9OkSo7bhdyfUN8Dq5QuksFiiuhJ
f1qFwuEPQjPkOuH/rlx6NqMTOsM3kzTUIwucvfG++h5OH/wF2nfeQMFLhy6PXeY3ra1/HPhPrlK4
MWZ26br+rYlyTSd0K0OxFiMgf77vEMhNEZAx9pkLky9tkWytoqfTJqYUT+v+clrMAfYPcqF04pvW
dGMd454cPd+vS3pZcfxQr6EwlDpmXGxr5PMG34L0pJgBe+0DpEni68zQDwWFUA1y/r+EkVzKLI/Y
1smW7Wp/NWQM2KmHwg+jqXnUTswLzJ5/5Nw6yqmooFpxp5VVCghgD0eGhwsOfhIV+qj9oUMdgve4
YNsVp4yeYmhiUmCKJWAnlh3uxuM69636/yE9lvw1To5lMlBcPIwddRIpnFyGTd1eT9zsVFzyW3Rj
+fTF/cp6ByG+pZQ8SOzE9rFTzKo92f7HEcCiKgy0cniwwXmNIasLslC0Oh1n0GUZpf41Jw2mNFFr
7kfDxneXG5U+goyV1jnrLfrOydGZ6YTna7GGiqnC2UP2O/gg4UKZnfO8kUflJruhdtgYKHCOSK87
LyrAyvR9BLWSfDFQrRsr9HeyrR04o6rznkZfyKrCrMR7F/U1RqIsGR+RNLopAX7VMGu1S7XJIPQC
TWY9UWIY7Doiv8eFthja5QA3q+mV+YnTcMhDqtLsremHoQfZOKDfPXoa5ZYZggkPdFwx76fPAX9+
lD8VbrcSBLp7T/XNlgtADQ9bd/nGOnQLMd0pMkIoolLaBpk4cACZ2SBwSKyiU4g81hAtOhAzcbUf
FdAAnSMcefLPIDS2aw4RMaMfkRkZH43RYISvontvyFKAOj1GcrneVB61/6Y8G1YfGKMKo94/1ESD
1fouBkUyoDJeuQINwreHV3Xqrx5x75SJKf9qVJQvTQKxNr5xBbbteb5VkUpsBgTpCYCRsuSUJxo/
hQPszWngsz+uV3acmGBLoX2Rgfvk74Nd67tIgkoiMjMZwEr2O6dv3LcJW6Wb6oDV2GxWQmbVfDbr
lZKbkCtdJC/tHahMmwHpU/p10IW4NPuYK6TZ3MCwCpIJS8HQLfObTNu/CwNIoSadvcMbSy48OpkU
36AY2QkHtcuPV3qP8LeBfrNjJS4NnP9dSaZnTG/Pc8G6CDLO7lc374enFeW0Y3hS5PU1oWtqYcTh
+CaDOOwprgmrz7NaIccxfuzcyPWenniBWXIsnxZzcSF2jK7gajEnOwfgcQ4S8aXHy8U7HIcHdq5/
/+bquBXJf+/pzc8h7HxWL5ORkMTzygYVY+b2boLVhaQXiX+ytGCFx+0YyJSOgUzQubGlEFwYYRed
hN1OvdzKDuBOPsoyYd/DqDf4X23fFkchdoZyJGUT06eI4gMv7jAd3Nq7im3tX/nCXL++DnKm7job
o42yBnDzdVoFFBcjlbvJDLOF3xIUS+Xmrzp2yPfW43fZCB9AdBF+9lnU0tV8v2gP7nNAqWbBTBCM
/t9+NgUcMSAqAYLKyDYhZcVliwNUuMxBXp8m/ms1NhO337MtTSyyJMddE5tppJDJJknaO8avfHh2
UXAQixBSy411nq9Vvb6VKh8q9Syjmx3rFOJw/FBiDcrXBe4XJbOERrNSuLuO3Z6HcIr9pxulV82y
cbnjwvG4y15jXKnOOCIImDOY7g1QtXmeFUpMse/3cE5b88E5MV9+3bwsjVJmfEz7LurvmNMF/fjz
c90NeIHw+N9yzBi1olnRC1hmuwbteueJP4gULnYBYJHoM8oZXjqMS4I29jiez6ZfS0sfRsazai3n
PkK/WVFUHt1X65vGIgGbztONxNzAsZkYctZuC7Gd40/UPK7BytVGDH9t8jhNzmRD1LfTMq9s4a12
JH9KK8uM6jSbWwMmpPv1OZITM/Qh+2PTEaa4YSyWie7ml/9bV4VLzeTGfwOord4ZFfzEAFj3O2S9
Jokb6m8wx6Peua67hTmh8QLv8UTXyu932XnkO0tGdHIs5Fb92qkUWRmczplhW8POLD8HxGte9JjT
pFMd5sDBkyIYspUKY7eUP06FmrE301dQ7OhDF3LmNw///0Ot7yg0A0SO3NidAqjFIAqKhhL4f5F/
q1Q+qRMsCcZ8hWYQR6T4sw6mfRih+jH+UdiD5/vXAErb7Gb9nrCnPantHP+2ieWXeA8ExPSYishp
HzW2Evx22S4J1c9TEqJXYBI4dCoVZnDvBPwuR85+wJwPurmIEUjFPKeSM+ME93e+2Xrb1jByjxwZ
xFnanDFzXLw6HdD3TOnL5MbHuFExjTvmv5OpHJJIXn8G9ScKEVOawjLSdQYYHTmPTVDp2j4O5DNm
mSWPFCq38jYFT/rs4FKYjQcEIIwSVgNI58kKnb2EdOVrrWhUdLaXMaziwKi/lG5Rba2laDkXWhD+
1ZPz8GBo56G2otP4KuKECCqvkDSlENbxBcljrXZDfoOSy3MMQlWG7liXKibsY+7LwdGRFmJIoZMH
7ZcnwCVSft58puDCBHOy7YB5YBH2wRDKbX8bEtLdNDNI7LEUYxSzsNOTTMs66x/vH9K9rfS7xqf1
CgHPvD93Q+b/TT/XYOzyzQQT0JGXl5GL0DI19MA44nzdg2a9c6IRTzD5CJg070q9e4vsLkdAqbKY
7davfoMIk5mkjc8jDKrphZao0nbQsGaAb8EAeTuvng3Cio3KJrGOCrJe7fVpPNb3f+ocZzlM7t28
JB94gMXVMzWouQ/h+9KtEG4N/Po98bWfzS419zpGJIySUhagR37/whxZ4CG9/Os28VLPuJpWhMmP
tSqhZ07N4EdhKSEUFfTXAKQrfdPdzFjn64LVdu+DZHpSs+D/6aXWC1mEaOOQ97ASBFiqPGksimGA
E3YVPac4KTCiAsNsr6U0h6Aqd93tYMV29hiIsAxD2JdhZBT4yzPGrGSK+2Is7lYGV0Jf7Z7Y36r7
qqC1imStCmni1pCfMLJo7Tx9RvlrbrDtWP1sHhPIzQ/MicHDemF/CHSHQJflDUXTxrO/Jku/NGid
HIMFZf9JPzjzvhIjrZ0KAQTXj8EChY3QTYTZC0xYMSz7BPSj0i5r8oWL4lCKx33NG0ENylA63N86
KCHV3AbWH7er4RICSUfxh2XHs97A15tK/KRCQpu/tIUcg23OfnF1H9PBcnOzLyeDu9U4jk3oT2/y
2hslm3e8THafp4FYWC7jG/tClpehMxAQrlEbsPJYLtWaRF5FObe1OagJoIuARgGa0QvVCBbiLjYa
ItwenBJCPdDjSYKbb12zbUTl/rUW3sWefYtqoG7Dkr8AK5m43Wb3S2y28OYidXj4oxtmFJ5pb2qD
vuSjUyxnw0+hK8UBoEbFkNVue9vb2vF+Bg8+ppMs3QpphKGNuRnp+YwQxiOQH15LBrIQzlDcg9fZ
0n4ruHxXBIHEy9kNc/o6d8F9ZCka6FLAPqkueK/1RUauj4x1zRzYBCctqGmOdUNZugKtJvGDZwdu
ha5IhBJlun7v3KUGTh2IWXqn5YEKHqsDpNlmLIn8WDrbWXZH0FbAMzMaCqBxNX7vUff4NQDLZcsl
4lgULiUhmzwf+FYeZj8Sz4G+JaZoiUq32K3xYrmkSubaKKdbR49DWGHW2pBFIPVRk/WjS3+Wy5dC
EDvByVYi8cDx1NC6G2/NTsExG0h2wBOQKGYRb6SnTBe5iI7pSvhQZYZcxn09d5GC5qYmLkPCYei4
t8wTYPFF7er3hg1d2pABYz9b6Kx8V380UgpgbldktjXYnGYbltZdttReAi4MzbOpFqVjyUVXMBbU
I1lLcQLSJPN968Ss6TjI4zCOg2FJgIQr2koBNm5QZEJ0F2sXfBDcw1Xp9N9WOuKgJ+cWOsHyzJxb
i9ezUtYd6jBZvEvfSfOk2CzMqlD8K/dCv0csyUS66aNuleVIy0crFUkjqCKEyjPvAaBjEd2B1DEB
yj7+xwXI5Kqmr3nRH6SpwYhBNwcCm4okDwJyP0+yQRKVzuib7CCEl9ZM2j3xLr8PKr7laj4RNzcP
tG0Yt2DNkGsV8oTAhu51Xnjnez4E2+hYWVNuQKdKRzQXHgTZbljbXLXnYEZmSOr+akUKUsxY9tP9
53ZMWbstXVSAkVbk13FxstyPxS9clslcnTlMQ/w40odH15k+3yC1NPpn3Hug/616HRhx9huzgpoG
RbmL5Yop1cl9Vx8zXYS+rHR7ut8PFgAeB7DAckInl+INiKYDmBfQ7M0AasfCVq7YnHu0n3gDvlLv
MNeqlk65YjSj2AJPfNybUQgZjeZy+vuXk0xvtPZB0Yk7nYHGVnLkFiz1wYQOficDiUITRdZqmUTc
kE1Hy/MVlnUDeNpq9WXwQN9TjpmYQrphHpJbyzgf1OAf1EQ6cwW7/HYA9FRQ+nF8k9weDWp2RvMJ
R6DDmqM5TBMH7npEAtKb6e3MPizUgy8+XZ9YFMz7c+NA0u72zPllqQPoj26Z6VVv2dBy73H4pTD6
o2KdhQOHnWEjx1e6NgNjR3oHRGR64/XKo2rr/oZPS/zJJ0h9iNy+CeQfUn8MgpDWOpQHiW46Xs+X
yRZDUOhS+CwCTsx8v+A09KXNu1EDwSnTPDN8p8JCFj83kJFKusOJuTlTBhZq3DTrxhSlB/Ohm60m
L4Bfo217g/eMeJrvMWrGUhXBQ+N0Q0CcO7O0LbJ2LK/BJkJRQ5nYbmTWqiYvwe6uyvX+/lmlEWZj
Q+ADT2NSyP7Pigjl6asD8PahHirhGT9LdKPTiZuYxD4gxWI3l2Zsk4xObL8W/Cgxj6YJT60Oxr7Y
4aDaBbK5QnvnQK2oWPUXX2BEiTaQ5CVqhNP64PFzog+wQESSIHXcjIi1ohop7yX4uiMK91X6Gn6O
8MltvnPJdFVQv++MHcvd/QpUgD4GFDnEHHVRBx5ibOIErtOdlmexpEUIHB2FgIMhYMp2/x/iCM6z
G17S2SfboWzlWD+juy8SZM0wPaj3HwCFoUweXo+TthUY7ZSu/mcDzwYMC5qhdDet02NZktrca7GV
dHWLB0pPFFXIzNFGd1HmPUMPmsNey3uBd5v87UQrgh49VBy3Xbmi6Kg2kt/3mS/EhDrdxPfUbLDe
H/vrpRFTPqkODpFL30a6jNKZqCQQKUUM8nrZNFXT8r9iQ1TGLdehoDEWWIDqfMtD0Mc5D9AoCk7f
i26MV6WDbDbRmVJa9LeOi6eg61BujciM0NSHsMFUeDnab6p51Rm+pYRJk/l7v3irkQMZ9qgm/CNv
BMJdHmZwgN1kh1wgExqhzTNOi++WdblWC52yRmXTj2YGy8BU/oxvTOFGrd7RzTf0vfzz0Iu1U0id
TNr35YMqhXr6x7NlvZJpUgydqudeR7UiccHqeP5G9h/sap5DgHqnxfw2OfFgETe1XNWwjNb5UsXU
ikr7LiUaoV0+cccdDq2RAAi3odWQcp+Rhj8OC1I8ahtc6dFqnp+nBZYGWNO0vaD+TtfbujPwlxbA
pb7cECtd/wH2gD1ary/MZX4jNoVSAe8acibP1CURh64SaIrh30PRPv5XnFXahEHoo1IMBfm9TcK5
Ddb87+yQn1w8L63sYyAVOh4azW2dUPBNIOEEXqrxdisyZkvpVb8Xb4apWz5egvcoDrW54m+4Pd17
WQCFrAoH+Odv0q4ImvXFl6QkR9qiPh51RNCHtTZty/WvF2J/iUo3m5uCObKhU//bKkpLClXETxBT
QXfHDLzzlnyNeh/s2he1mvJA+sDMFZhXm4U/Y03WzfO6QBZKYT4VdHT/Us5B500dISCl+6qbWQXX
A6Xp5/f8WJslattX6lVVnVI3xvz/AQxaoQlxP42MVGA8mcdK1sdKnoDsOp62CjCZr1J/EqMTAfgx
w+8mptt1WnW4t+GHta24nw0Ig2SXLv8GE1OxsE8XeDRi/2XmxMF5ZN2mRXX1B9tZCZuuxoYXUFK8
Y6IHIIZcdBnwjnH12VsKuNi+OjLKpZ6LNqP84yeqL3gNbARE3yIFpoV0GUONtCQTGT5idIYnaiyG
jyfwyIsqzJ5hra2NvjQNxU0k+eU4gjmSTPamDTznZHoVSmCvMxYXSkCCCdoVPpDFDVdLPqImuKcW
K0lJ+eCkQcecmIkzjok20rrH6qPOeL68Xbccd0wrR+l22vQxe9YWbW8EZ7rBuBteRU25wIPsbB5q
MCBZeDbeQjN95xofjxd6Va0pWc2S3cGFtN6NU8+udvQBYOM/6oQYMpQvWDxFNg1PajkNq9MBAok5
gBPEhFiZ30uuY7bVXyCIczvLchVPdsePfXYv9mu1FhFBwmiVyS2+LGa7exR1utp5Rhxt0+gYGd8a
guedf01HZw7eCG+YflAekU3gqTwl3dr/lkBMg0HXgJN9sdzhq2ct/dqKz0wVqrkvaYpupCTZJDJo
lmVfAgZa2ks3/khl/+GfxQQmx5kRzGGanwZh1BJYrK8FgSJ7SC0EhofoJLVpLhHtH8Ow2W8USZVc
ohp3MaB0cm+S78lDX1aZJdeyDBryJDlnGHaUtaGuKNW2b+khXa7HPLhRqD47C4e0K1PTYjrWBB08
oj0kMSSEH8zLkkZPzBRGnn4NZ1fJLFUW4oFrQYQUGU31EbEZjpbBW9/PivIIQY2DvPU7baLR9zRq
gPoUMXqlTzRvG50kSZI4si2nxW65Kz/uS+W9HUo4B4uiQ8wg2r/EaBYVEmFBfO+eHHvCapnwW7+G
jFj+Z3346/bzJvNZNoW2zHHLAFPqQkzFR0BcFjhBfBhDNbFowts7iKmH6cysrQH34Y6eSgtcLvHK
ovBNEoT1Dp2R7bO8T8cHQeowzcgnHN004C4KP39s0VbMh7aQ7q5sNvcJRj9gkmcxMRn5Cit+BsWS
3hr9gXgxwxhf2vVndYlgL/4T+Y1/dgfh8UaYB6bZwmqaK1yA43/GDyjpC4syLy5llObcMHkBvyB1
AdDLxjmsqeOvwoWhvlvgt3qlxGus2BNua7mxBuBw8QFwF+9xHBz/tGHKyYvvpNR18w2uPEyMZ7ns
WcQtOWMq6KmOHDLFWErn5OZpOyfHmOITzAgDr362/DhrYEOwRthDnwVBgE12/P0Gcbbn/kB/jCn9
L2INCjrVqypNM/ItfN5m0LafpOIzLLw9BXin9Gf5bNhr5FGJ//2V8C4QJ+6QFAKEWyIbyZO10aUL
AT8he2Kx3bcQ6a6JnI3IqFbi5QT5goi/JCL0+e9kU3OBhjHYFImT64sf/lgDK2iQj21UjkaiKOmX
DMRYm1Dh/FmeXElk4BOr4vRYhM2lEyGL0UB+D6tLjWLiRGAHBR0NMAmq8dp1UNV/a9RlRIRlmIOc
KqwmfYizc6UCegHNNB/UHD38jFbDU7WgbQIgutbJLOkKuIZrwFzxz6TNQxlDuA21XibWHMaCzF82
r1h7+h9LU8izb03hjaLjuDVUUHASf+GFr3uzD20lTq+Zfnbkmef7D61EsCnP8FaFNYnzNMpa7/oZ
Eqt9PC1qBel9webkdXA1mav2NoXm2sNm1h/O+FSS9AffZ9XgOGQN8LaEdUlmjKGC0pLf8nCrIc1q
imCiV8eDxZkSjYgZ7gIlemVm4YlIJ9UIjSYOFD2/QUzfVvfbCGZ7HTSsqlApUycDZ18nPxjytVI1
OdHq57b2BdGxyGZemRqZq5xbb8XxzHK8aJq2wPEy1rjIwR7+LMTc2ZsCdAxOPw7IHrH8D0ZgvML+
pNq1GKoooQV0aOY2ZYacspmKhbz2XmHoxgIV8R13l6gHeOgCDQnM/SbHzrUd+JDhpbsg/sVRfEZG
qYvpd8xMbBpukAiXC7IKmxz5CyHSC5yFT/UX5ipc3bJiT650Sn4uSG5OL9G2YxDDsw8c456SDiLL
Hy0zZcRur+GjvhvmJVqCevoXUhnc0hmq13pA0VFu9VsNgYKm79+xjVvMFwurFPJIsy6+6eDggUJO
wA93g4p0WRjsgq2XO02ktSL0SrrdB4rRZDaj1NYN1HO+SAzvDFHTnpTXV8ElPewyqjWMkKegS6lj
lwpHSJ8DcCtNlKDJd8nSgDrZqAbMHDwF30eky+xRoAAvYPCxxxeKa87kTRTlNCDRLc+ucQxtyWhv
uQyc07NeEcw4RZnQdtCovRWEyIruVj3AmfC0B6JddG0x6/lTFYvi5eP7sJ3Jr9am86NjEyF2Hc9d
d9rNuAgClq8ZKqyLzUkJM2y7+L38XKVy4DZdV3l55GmG3zQlBCOntyvJAAGX1Nh5W1krqzlv1Bhg
ERDG+r/sayD1sW9nVEoNvs+xq+HrQfu5v/IRX0tVVaw23+W64my5Fxp5e6YtQvTPXth5ivFgqHc4
253nxjRfbw8pw6foMOPpHWt6Oujf4XftlQ5fV9CCQhFp2Aq0QgQST9flfGguqNyxpgUxvnd0qa4a
5eyqVeVxQdNEd4wRv/LVPcGa1gQuOjF3RJ1y6RvUzy58Qo79aIByOgWKRL12pTIpMIigp0/nneaQ
/Z7vgmLYW95HBu9lCnRNwmuXHUOlgboyid0t/Vl6eWOyHon/7iFQqWTdEKknlQX51Xp4IeKumNZQ
P14GddKwhdFpplX4GM1KNk4TUGD90QmLmayxCnbfbpbsWQzO6TS27M0waDwcxTcgR2xiJte2xKJ0
cxf+r5GxksCXPt2mEXbGAf4nhZMgtNM65GECjrUuRxV0S6ychQ0QXqQolz/59J/Tf9I2jJUPMpy9
Vum7O469t142sn2IrP+nJrfhj5ECH4VoE7CEvlUjDW35mZiNLwPVHQyln7LlFr8gE9EYiEdD4MFo
PGVFu2F4oL5PGv6CZQjn5O33rQtIqDYRZc/vQ5BEzwPWMcMN6uud6+s0QLQ85mcdebPA7cQ7C4jS
7Lr3kVJTZxsc6pUz8NV9OO9otex22VPPYzt9N1Gg8i4yQDJDncajY/oFKqSjgAoh9OVZKt5XPM/Y
JR8Dt2Xq8IHI4SZ6UTco9WOtSjZnXv/zOS/qMoYzVhJTztCxbmGzI3pbjxQSlFx6vmBFrxtBFyQg
9T5sINmN9t/sw5kZKfbhdMzg8nLeiRG6aIelDPMcA/LBaWG0SZ6QeYgD9JN0NNqlwz/QwOr9d4Fo
5ayaoqA6uz4tZThKEp8nI08VhMDfDxKjKY3Cfo19AUoL5LJdeX4+xlx/j8GMtv0/mBo32T9RGxqy
QnoJQMbf/4COMrAOTopFv+G0gE07ObyvBYFOaekgu5KvPEwqbelYuyaiGvi+TPH1dG4Z6ENvrAxy
JxjfAQxwmkyeFA87p3NcDOLaE+7wo/kdDKi2lO0WLRNZMiEGxzMyeatByXlVlwLrckqBi00j2hBa
UJ5/cvyhVYnDdDO0l0uzo3sniaMhJldY9i+bOBDhC7aceYsa6uE0nlPgMZKC9VyDAS/YNDkd8A46
iBCUzYfErrZndF9XQl/eJkYAItCXVAOBGJFbSyUSXSwUaBp4AjrSv4qlqXkWLcRGL+ehUU0OW1ye
vhs7O143zSPrHOrgEfBbvb7Eh9xuBtLneo0LmGuId+EaZpK7burMN6W9KVjT+ZnoAFMBB+9+XjoP
CKgoJufBSWMUHTcxSKMKvlw46jVnPQHAXCdxnD3mY76uY1NKNzaCW/YLKmuRoURKgbvqvehnUlIx
C6jJiVNGmCvdXca2/Fn/w6mI0YoIns+aPpFkPY5ej1tQUVXPDC/JFBlpymeisK4o6UcKeN7ljZJN
dBD1fPt+bSvk2Q/Sl36bt2GRzRqYIVejY4i+nSCFjh79GvvrvWZR+sF5UFNpNqfUy73LQoDgI872
nBTVeQNcRIizciIEj4EiJPze3FPfo/o8lrw5odSYbNOmjqNig2PXl0HZwcmUpoHWaENphmBKFGDe
96Sdt6Y5B/f+kVJWIYjTyyc6lb1LlFGOV0OruWR19qLSTiJObl80oSpXZcBXUIh2E2qL+q1LQ8IU
56xNZaiKilK7GUgUIbaVG51dK1hGBJtFXhILfhHtYVJeYRDy+EpUfKaNq0yT8AVwNltKtcdRFSOG
OPFfs4z8SogvixB4jDE2aGaX0urX87hrHoFxx2dzVnxWSnD/AnT6z37owzv6BZi2Uv2AwStQbrul
XDXckIFlOUGtPZH4YHf/bSTDAVj97pIqzPJc5JZn7wf5pWBiCXFnC5eH1THnLCHfJq44sah97n3I
8db5tm1wONBehuN9G5IEoLHk2pm1tKMaelhKNneoFKjBh7UN1jI0btfnl0BjkHOB4jCj1EN3FK5g
M8o7tlce1hb1gBbBfYhsS5Tn295nLVrODV1In2UKyQpw7TBHHOIjdsJ8M6KYPK3y5uYB44dN8UMT
KNtdm6FyRnppkICpJxfCn0k+7opwuuYEivwaSUz/2RCZRTnlwahlBJjaGd0+AK0YKDkttzJ2elQz
sZGKasYndiD8zYNOJ3MSTH144uT2t6KXmtAP8FixNqNWYAAKhKWwIngyCJY4w1UYpHIrYmn8fJUd
YhOIm6Fx2X4UnlHYBYYTjLxtshxGU+YRRwuEGkamXsDVcKL2W6hkEHVCv0ZW3/HLvoYqNo8gKJwg
YIWJVVoJrJACKev3laYmm4HSvG+cDEkCjCT1ChQNGhM8948cUQ7c56wGCm8ztiBP9kIQmjm72juS
BVvEZqgbrC8CEF4TiXwMuSe43pmaUu+LPEYlLH9nlbSb1pOdazCVzGYQFWPoniYf7Q3wFPbOrfFj
PpwVGaW54oHkU4uvKNNXnlCiOVimdv3wyMIMaROfZGrnyU3LMBHHobHU+/pSa7I4mhwaqapdxTcP
KIuz3R2rRQAZCzDcYuRK9b1YL6Y7fbWsY8WU+FhyqEQfOp5Q1xruKPk0IXjdnrbjIRxY9CNDHx0Q
5g/vxq9s6rcRJK1zT7W+urMlYJbpHDL7
`protect end_protected
