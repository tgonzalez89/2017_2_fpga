��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR���[{�T���CK��TC,���:�
&��d!��]9�'D`�"9 S%�aQ�`!�6������V�W�l�a锦E(�\gC�slu�4U5=1�N�m��l�9ў��P���B�@+yg��=�}|֦���ָJޒdm�^��+��d)%����r�&���CI�m���֜�H��y�>��Dד9��i�5�^�%�"i��G��B"��%Kό�a`#,jb��!��*��In�T�*����:Ib�����]�e��K(�&x�;?iX��pٽ��I����=���Dk¤��4:s;w��SP.A���邼��;,o\�N�"T"m�:F��,BC�ۃ=zC3�5���@����T�Դg(q3�J�߶ԛ�ҫ-1b!�
�����Ep��L�X6� ��U��l@���淟f�_�}Ԯ�\��>f-�3�D�lNw�*���f�!}9F�� f�^���ɛ\�|Ƈ������s�p*�Ƒ�2p♕��,��]W��.���0��3{(	�4^��'�/��ÙV�g��"�	�@�PX����󔞫��W����� �B�����I"�z��S�Wk��o� � ��g(�C���#+�Hy�C�!S��	��/�J�V�t� ���*V)��"���fתW (H���j�S=�L�zwkj��ҏ1N;��5PL���=o�-�y�ҿ�^��m�'����c�IH�{ �a/*7(��7׫H2a# h�z��I�s�z����:|¨k$��W��4-��a?u�o�쁀�}1�^ic��L �WiHG�@ٸ��'L��MD��7�� �{O㾣��x�������-�S�bg1,vV�� ���k�2I]{(&ʂtj3k��`]!��iV����݁�8��&;F-8��[���4�n0���:���cnUo+��!�Ia�`��&��ՙ�HY��o�;�A=�p����i����D���~l�p��l�T>��nw����I�E��w0z�U���de�V0��Њ'F���Sw�0�EMtjR������^@w8�_s����c;o���0��m4����x�I�ei�_D���e{z�mx�Z���$���GG&������8R�`��)���{-�6�dpi�K��ʋ�����^On�v�ww
Z�y�&ʠ�ی/�4r���'�>�ƻ��>��΁s�R�rv�Y���ٴl�޿��j�
#�4�=�2��N�C�h�hE�����3ޖP��u�I��<��19�!0������@ϱ#k��#~8M�U�`˴!j�=P��IM�D[l6�ЧH��we�9Jy(�PBͦ��p�)�1�T0�����6[K�[�P�yH��yzN.W��)Gw�Mt���?fx���OڥIF���p���Q�����ߺmV�"�?Շ�++U�l�� �i�T�q���A,���d�����FCn`z�՗M$�z�*�u�p�ݞ��naFg{� ��P��Q��i�[�ōI�#z�Ș�/��+4(B@S=�ɯ�E#��$�?�<��"T�>,qѱ=����6c�B���eu��}��r��C�4��qAu��y"%�Y�0;@_�E^��%h�.u/��_#A���Lz���<w�|6ޗ#"��f����P�s���W��c"����R~l�#��#D��S=�ce2VcM���"��е��w���P���_xAiFGQP��)�ä��YH�W��*2P��"V�1̮"��5@�������nvF#v2(=%�����N�C���ɧ�kj��4�f���t���X��(8�TP �11ڧgӥ>1�)tbtp5���8t��A����ˣ�oS��4߃��#d7ҹ����=�~�YoD+eMQr��\j�%���Z�������4jzP�����?�o�Ѿ��[�QX19�V�A��	������N��!�2��(3�a�`�:D�li)�-�-���xFX0��m�A��b}woM�ZK��|m��|d7�6�ۉ��}�~�G�:�����(�69�J �^51��0��^�)��OC,�J��P��܆
��}��T�,��e<�.`P���(�@�s����E��wpE�4Ǜ��/"�`ަQ�5Д�M���>Bh�z�1�(��̈�� �;Q/�UN���uL^��U�TԦ"j���1�PT��dF��.�L��7�d�4ڸgHX	&:/,��S��iҞ�1�����
�Aҕ#|�^���NS����W��
�6���c�hT�_��1�-�(���Ų\T���Z��q-CN%���̶���*���4j�+�+Ff�eI\�#�D!��dB��jG�?����σ6���b��x���Xf����P%��q��S��r-#���F�?�������+�e�ߓ�A�����1�П܈9Ӛ����&�ݻɕl�tAZ4
Y���b|~@5Y��_#�Q���ǆ��$gy�c��׌w�v��s)�:�dL��x5�:�=���	K�}�y����)��JO[���j�ݲLJ!_���R�.���y���M-[ ���6�mB���Z �`�/P��S����9������j VpN�~���S�Q7�3.$��w{B��dF3�I�$�J[���4cCzq��+�j�$� ��ޠ�xD6:\o�I�hi�ΰ�]�C�JT��>� �rq�������	�Љ���˗����Xo��\�;�Q@xNG�N��T%���@f�u팻��r�8��#���?��d]�T�r��kq��Ms/gя����2��ϖ�,�:fe������jp���/���3���"saz���&�&�1P-0Ns��	>Q��q�>PAՂKaQ�
dsOǧ�����ub�P4��^�O��U���Hk�T*:��L�sɍ�C3�����Y]��&@!*��}�/�P�GS1{?m�o �(�jJ��_Pf����r����#f�:���o9hփ�{�?o8׸|w�uo%J'>�1�<����^���!�#�e�NR �.�:���uO1L
��׭�Ė�P�7��1����*�� OwLe�]R��,P��w����~�Q�ʧs�9��:r9w��l����'I\
XU�F����9� �̕C�/HO^���R7����z
p��tl��T�d�����Y���N���S]��v�/�>e��&l��f{���!ʰ~���F�3ˡŸp���πk���W@<l0����ͭҡ^��>�A�Q��͓�X��P���#�U(I�-�L���Q �����������@�����b64����uL��G��^��F�"כ=3]nf��siڎ��Ҋʧ����,U	Ʃ8ƹ����f-nV�_4KFx�@U�4�f�����mv_WFi����M�<L�^ %����+�9ލ�E��j���9��D���_�S��h�l���Ғ~�dt����Zb�3S7�!�Cs�G �2�v���D�0�/p4"C���/�v�^��{�b�v�dLLWU�j�Ґ�S��L�뻾Uoڒ�&{:�b�� .��]_R�^'h\G�ORbuO�q��?���� ��r��x\�#Z)$^�3�~(���^�"�cqK(0��"���`�������������s�u?�k�>s���^D�����7�5��8�.�riPK�X΃�x���HHؗ�O���>nV{6�8���m|W�ء����ƙ-���f���!��U3��ȸ�����<��e�k\)*޽N��m��nq!��_�O#j�o&��'���