��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR���[{�T���CK��TC,���:�
&��d!��]9�'D`�"9 S%�aQ�`!�6������V�W�l�a锦E(�\gC�slu�4U5=1�N�m��l�9ў��P���B�@+yg��=�}|֦���ָJ.�&L����:(?�6Я��W�j��5螈������p�2��`����(P�k1.y<��p-��kZYU���\/���󚇖��2�t�O��6T@�l8xN)QӂM���ԩ�N���8�ZE~��.�yQT?�i��k��-�T��f�ڑ7W=ם"(�$�EW�"�[��C_��{l����T�C �xw�}���,��JV�iU�Jن����PAB]נ��������\`D *�^��P����e�8�;�5>��:��x��������L]Ї��O�����K>��r��摪R=s�`�s}U� wU�B�mM�2JC�-��tW{m? Ӯ�/�y�!)r�� �p|�Wu�ӻ�.kΌ�g����d��h�%��$1�Y�����Hk*	0�����9�[g�s���4�n		3��z�"״�ӥ�1߅3�9���j.b9�!>�F�䓜�M��W��Z�j�����E᪘�ր�}�O���^Iw�+cA��lq�,�z(�-�y�i=��P��ZS�F[d����af!���8����`��,qwe��W�L)ݜ�Ǘ��k~x�9=�C�/+͈	��SB�*��A� �n�}�sF�d�⪒�jh�&��\�����U�ݿ�Z��U�b�����h(GDUV��#�DCr������[���+YYZ�\�ӋXi囨�a�5�]�G��隮!���J�S�ѯR����/r��ng���
Zr���/�u�N7. ��
x�{#d#���	:��W �$`r����.������(O�[go��n9mܜ>������.�c"��i�B�-���N!d��O���n�����<�sb6�%5�*��D�]����w����)#�1PV>�;Y{���Ja{0 � �:Jxu�͡���w�p	@rX����.��F��wi��$3$���֖ѳ���>�>���h�<imU�K�|<t�e�]�QY)��~�J���������*�A�����̈�2B��\���D%�w��ApgF
H��P�H���tB�\��]P�O�L��Gv���m���D��@]r�ir��=Ʊ��q���Mǳ�5�dFS:�����r�RlY�X#&J	�Gm�L����F�2�C�8j��c�ȥrȗ�K��e�����
�0&�D#��7
D����5��k�� ����}�!��[Mp�=.����uW��μ՗?ܼ1�v����fU�����pG�T��_g�e��O��s��*�{5�%�P�$Q2n�]�>ES���ؿ��8�Ka���Pw3��N�z����0����e�I��r�4�ŏ�ܜ���
n�H��J;	�!eV;�-uM�����#�tEց�\Ow]�@��'J�RB]�g��@�ʐ��<d$���HJ��8D��,����S� �|fۖg�L
k��l�)@5��
�¬��l^z|�����߯�Qd;TKO	�[j��)\+�1^��TM}M~c!����[��i%�$�,3(&����������#���Z� P��X��S�����.:����SM�jV��q���v諛�3h���DY������	v�'O���x2|≥Ȃ��d���R{LQJۜ(�Jz�����}t	,���M`��:�Wz_ �{'R>��a�6���	���q�H-3G�/��=��6�F2��*T,cF�Ǆ˒qG������t����]&8�q�r���[�WZ�  _w�00�)}�����p�5{���Fy7xyo %��Z���\�n�?��.b�'	�vaf"�z���@��V�3z�|r%�;a�{���(t޿ ��UK(��M��0�H;�+WB��T�������;���Q���F�H�3�By�o`���K�S1��kؕ�:��Qf����V�s�=v�b�E$�OF;zM��4�͡y��:"���|�B��=��w�Dπ�~	!n���J���P^盭�KY�w�Q�w�����_�{��xNܿ��P~��'`K�|�G�L������)4xLD�4��.���os�=S���ըtD3B±��a����y�Z�ZCn����.��3���`���9����m�r�-Fᾓ��r�-.]	"�:���s}��>Q�5-�_ dL����'�[��:>ݮ�§��h���NY��ɿ�o8޹B�Ȣ썛Bq�u@���f�Ǯ2��v���������C'IJ�U*����7�����ۍdbA�"�G�^����o&�'C� ��N-Y_K��`ݩ7%��'W7�x��������eq���P �M�k�EBS�Yا{�r�)("fq&++4@��7η�2��@P�o����K�&�^��=�(!�_]W���Ahg��.���O��̍�Ϡ΅��?�N����3�a�%L
f��oGro���v�/�or��F�����սHD��5F��;t�z���>��3�M>�ff31�"��>��:^v�|(��.��2t���zrm�}�N�������_�v��<N�y�|�+J���Z��r|�R�g�}���@CD.9���ge
���W�$�u�W�q�E�x�p�q��gҦ,�׊�M1�x��>�tO%u�X�g�%왝�6�f��|Q�c�SL a�J���� ���mQPH�*��=��o��h&Nݨ�©�\[�;�Σ�Y�b���|�#ћ�yZ��ߖ�lf���̙H�h{
������,�Rf'xo���|�^���$��d5Gi�<xh��Ƞ�=t0%F|p���nneX����X�M��o3�%�W/�]IG��NMp0A��ӷ&l�+i��*����bU�Qq�{�>���:��9�0������M��ʉJb-�g3��ǃ�!>t_��f)���	��7�WO'	&0�� [X�9hN�O [���][�R�V�-~�iCZ[)��#p���P���R ��<��gQ� Y.~�@Ϛ*֬<����qH��|}E��r@���<���c"��o�7_hv�
D���b9ϑk�b�����b�i�I�6���wB�*ND$�U�k�StR=UO*/�9^aBO�zUb���P2�]
3hM|Z�*�vhb��&�Q,�Dդ�q���\���ʡQ�������|��9[o�U`��:׫Ľ8�����N�ͫ3��8Kf�t��*����{c��-����.a�=�k������mّy��l!i.:��^a�8�NP����� ��d۷��vW*��˓�^�����oY�a�}��y�}�\��L�]
��7/��������9���G��(��R%�ʎ{G��?.��szW�r��.��4�S{4~�����|�|_�� ��«��d�$�����c�:�&��:r+�|U�ؐ��ьv�k�;X�PCW�Mj���ك�޶��'cX4l��43xa�>I���Ǹ��
����{@a#����f=����r�k_�kT>H�$����˅���/�$�O��|HX��B�6�_�NX�&����H��m�Z���#�P���醊U�Y�կx�d����Ȯ�]-ה�N���5�ö�ḭ~<�N���6������n?j#Y%�����s�+��*��C�~E��b���ziP�q%3#����&]�<�e�޸35�w�>E/!����/���N&�VW�١&�@�r�M}���id��]���g� '�d7�!<�-[pG�ӿ���/��+t+�_qSH]-.�.�-�LP/_��#��x%�C#	�M��a�[H!�v
���ʪ�h�r{�2��l�^;j�~���+�ʈ�3?L��D3a�������L����ʜ%�ӹq�qR5 �o�g�˝|�Y�ߡ�3���W:@^���=���崖����A���Yu�T��*P�>�`�d����k��R��b|@Dڟz�N��/��K ��sCh����I@�swP;.�Y䒲:�3�h-߀�@WS��Oؤ�C�c��~x��)�$�!��c�Q^���65���40�ʻ�.0u�eb�28F��_�zZp���$�J��_�l��.��{IR{{Ch>���u�FOlq�S�[�:���}s�-�E
u*�\�
qO�[2���	M���9i�x����`r����\~�O����
�3�eTuS�|id�G�������ِh��[�gJ�6�nԹ(�쮹�f����u:�۔��� ��$�jE?�Hea)�j�zR��d�t`��
����E>��Fa�HP��`u��U�up�g�?`9NqzUb'�Bm�+�mMT���^\9�#@�қq�m�@�N0����Cu����L�Gv�=����<L���X�]��
XvB4�=Yh��05-Ս2���F	� ]��|j.��[��}Ä�G��1�.���!k��&�����F4�SZ1�v�j��΂��h��H���e���ٴ�Px9�	��2<�����1`��W$^eҷf-�m�ˑH�7�}9���ipo_�ӔqU���y^鞈��)�_n	!��4��XU�{;#���(gq�Q9��@5�m���q��O��3�Y����[�Դ}���,0S�oݴs�E���_����z��{�R�D����KW�<_5�#��6������	*G��=��=���fN��S����E;�{E��c��T�V4�a`�';yl��+�����l/��r��c?3�C�:��f�j�K�ߨi�۷��bbO݉'���`�=�W*slV3v|Ww�3 ���
P�;�� W�P8B�7EKiQ�r�G��}��Ih���X8ǔA���b��_��4ۚ�%���`�k�$�W~�mE\�A�K���O�{����uECNU6R�ز�a������9qX���KV-��1/����3���CS��E�F��Tw7�x�X��t9xH��%ކ�.����J�;h�/m�N���s�+��i�����nʊJ�.��#
Z���GJUӂ^z
q��@~����r�	��r)�%��%Hz
���P����Tn���ĮR�B�NAf��'Qd5,��@Y�r"�h	S�r��Eؒ�so�A�T]��g��5[KZ9�P<�;�٧E�7�̱���'	��[>�	��Z����wp�BЛ�9�Ť�	��ZU��pv8`�p2�9��G���xǭ_ҙ�|d�q�䂥3mf��;B�%ՠ�$��*������qq��X���Q��e�܌�󎅛5�^�Q.���"a���$��y�0iC�'uŭ'���k� �_�X
@��{�C���DHL�k�ڟm�M�e#��r�YQ�p�7�㳃$��xe(�����2�mo��$�	���շ)��́\a]A<��?��gGF^�ؗ�Ư}�[��Ӂ��\x�$�G�7��%�ʆH_���os���=[$� d���p^��"����)1��n�.*t'b!m�XK�i�˯򀜁�,�p�Z�;ݘ:���-[4d��@���}����2&�jv�J�l� n?���Z�V��7�J��s��F;�0q������gI�b�;��В��p�a�֔Ѥ�����AN][�/c��쒿����}7R������o#W�Kv���p�w��5j���
�Fo���72�&�z�kJ���\4.�{�Yf��B�5�\3>����ˇ)�-�R�5&�2{���ߠ�~��j]�ǴNt<�5O]6�>�*����5���3y�W���?PY��W��9�9���I�;>���|�k��,E�%�]Q �B)}��#-�[��=7 Ml+�QQ��mP;�T[�P*���j��f&�������B�S�߲#ƾ�<���7F`q_w��kOb��)#l�:��9�F۴<Yp��<�g3"9b����<�Ոu�Z��أcI��kW�WT��zELn�C��9���­�T,ry�#}�"^�u��B���W�ؕ[�u���0I ���M�YG!:F66�=T� 卛_ ��U�7��J�OQ��g�q�R�*c5��>B`�[��s��P���X}��^�z�=������]U����mB�qB���n[�KP���vGAA��VDЇr`n~�z�@/덮�³��k���p숣�(�	���?T�=g��&�� L���
aGl��H~�f�)S8��s������f�W4O��OϘtT��-��3׫�s#��3Ҿ�|0"�?�����#
jo�������D'4��F�I.�P��P礥�1�B�[���4���P,�Em�>o���(�٘.�0�ګZ�;������>�6���=W���
����$�J*�M��!���.ľ�V:�l�s�l`
�
4E
���;�q���_U�=�-i�d)�{+�֕�l���=2�p���(y#b���?<��8�x+���{�\:R�͈Mj����'[{�����z��?��<����^�|�M]!��z� �|a���"�h����w�]|�3~�ʝ�{3��9��ƞ�fo�z�^C+���)G���.�`�R�Z�l�a�y��p���x�h���h�,�
gW�N($R�&5���)�w
���Yػ�}�"��q9bs�h�[�Da�W�8��Akz���)����J��v�N�a���H����^��6*%�#V���D�u-m���G�S�,<#���O�,<�h��-��kO�:�"I.��^!��U�H�>�>q}#B3�O�mӶNjZ?LS���VkS�o./�ک�W�m��0� @׍��w'^��^��1�<�xϪά��q,�aQ�k5r�Od�gj�
j��y�2V��?�4����(v_�pr���&��|Jm�!��+ٻd�v>zb���Q�ː$����.<ux�mw�h��3��v�`7�ՑhRR�i��?F���1�z���`��� PB-�Q�P�DSY �˹�,)'e��M!��?T'F��ҭܯ��13*1L�ܒ��:����(1���:j��U�v��~�"A�16�bw��|��લ��e3l��]Vd!�=���	<��p��v��U�‎H��z�7�����5:�kz�����#q72�^��i��N���wʄ7j���%��`�1.����q�|Т�^���SF�)�	�A��Kq+�F�Ō��(S0I����էƘT��إ:���
ۄTmr�l���ؤZ-i�Vf�.֞/�"~�B�v�&Q����s��{&I�ݞ)��2>I�$���� TФY/�V�+��q�b�jd����C/�@S�]�ڏ��[��I��)+�
ed�w�z��F#E UEN�ɥ�laRÁ��S���|^�M�q5y��KהcW��"�)C���6��m�Y�8,�͊���`ΈGH��@�ǻ؇]Z�L���,��4[ko��(+67�(��6�r�c�X��X3R�k2��	�O
��Z���Gӣyh���>�|��e�#��6']�e ^��ͨO�z8r�sxexgJ��\�Le�}�N�������s��G�m������#6����X�[���9���h$�f=Z��[ތ�#-�p�Qu��Z��H�WjX�N~���Z	���#�Iwl��|K1��,��e��s���gY��V7�^U����I��ز���N��`𡒺�1��oRq^���Ѐ@�i����9��JK���xR��nb?a3�z��q��q�؞ǌ&�l���U�D�g1���U�M��K!8|��7�u�ea j]Y��w�%M�s�r����uܾ��w��w�7pQf�7�V���\ ^�=pǩ��:�39t�h��
�s�S,�^`�W�p�?pzvx
(Oj��)��̾��
Du�pGH�
IӐӠ�-��;�>�`--!�5Z���4-�K�㏬/p��nM���3�@Tk�?E�B*��>��
���mc+�q���`)'��l�%^?d�o�[���ڋ� t���:��C���C6�-�<��o4��~2�+����dh%�c�+�B�����Rf���Zs �l�g *���l��K��#J�hz�e�Թ������o�=�4[e�rQ�H@��ő�8Db�T�����y~��ӝ�4A� ���+7#}�OW	w΋���|�@�2�	�g���v!�7�R�@ɼl�Q1���:(�(����#q���K�k���>\��+P��ҿ�8�f�I��e0ī>�P	}���K�Z�J�#���֕�#��)�{����;Zve46��HR��G�i�Qu�֧9�X�(*o@v�s���u�/��6%!��V+��^`�gbyW��<�8���f�� g"��FYM� ֈ�z��?ն��W��)�]�iA{�߸P�[$$�2"_��E��7����Y�u	Im�jZ�B����M�j�K��O5�壭a�{��J�<(7�HZ�r�z%P�%�.���5��Nu�]�fA☟��&����;�+z5���<"��Z%o��F���"��ws�^��	�ߏ�t���l��\6:ʐ���/r~&���U9�h�J'wL��}�Ğ� ��5�gn[���ې~��e��FgT�����Q�4�b@�b�b��?�r�S�����Z
�2��g"��ݑ�h&M&v����R)��#ߓ0���jrb�x�=E!���;uOSp����5�i3z*�������}�Z�5S�g-���3ōI(�2L�I�"*����P��,��T폴$�b�{ �hF�|�0�ֶU.�R�(G��l�'�8B����qM�p� �eؕ��Sh���}�J)?�)������P�����4��U��O���cR�65�Q�1��1鑴p��+����U����!��M�
���#້$;ҙ�!�i���fUˋ����Zwc:��̇2�H5~��2��q���	�4�\�N[����"��յ�Et�A8eܯi����"A|'���ރЉ`t�����aW��j=�G�<";�h3��٨M����1ϰ�U%��܁�����˕jf�d�G�ir��33␨ޤ�f���SE�Tǉ�!�lT�mԻ�n�X���߼���|�`����{۞�DP�X�"+�'6�0�ƾL�LK��C����?Ʈ
S6�3d�!��50�m�`'�u�"�G�u�7�-kf�?G�	���<-G�;%��0F��c���9��"��~�n:hF����7u�%A�=OR\g��L�v�I=�^�َ�m��Ł�~�|/�q���n��@a�#Et�rt�8�4�(��ɢ��HJo�q>���+E&<`G]x��k�S��ͮ?s���Q�щ�!���C,���"#W�r�9��^�q$:v����J��WUkm�-���@�{�(�NgE�dx��#���96�/���9$�,�
c���-��K�.���\O�j��)�$ss����ܲ����aJ7
���([C�=��߹1�wU&a���e­"���31��S4��d� ����V����y��I�7����x[��e{�|)��]���\V�����B1��8w�R����/���a�>�}�FB��Z}���V��^-f�������b��_�Y��o�5�MG/��#`cm:pq?;ǘ9a`�E��pB���ˬ�T��m�L�. ���׿�x�B���@���]��&R�ԛh�p(EQ2�!��B{ٹot����W;�������Y���`�~eK��� �r1�$=u͔�李�8�K6�  ���i��>r;L�<�s%� ��6�~nh���*��.�.�u��B}�Ƶ+����U�"R��2�Ls %�Mx����!qY�u�i��5},��o�)k��V[�]�èF� ��D�y��3&������ﶈ��bd�q����{U
N��&���-�zZ�e�s��<�^��%� '��0�-f+���)k�麏���'u��H�;�B}�
�Y�u�`f0Ĳ-��ߣ�x�z��##�,�+���H4�}�����c���epQ$�J�%���E������<t+E��]��Y��B\z��p�M����P�Z� �ױc����a=_������ھI��'ص��F�g3���gV�����pM��[25K����P����/���ﱻ�a>~1�eQ����V�J�h��:����k��Ƅ��㢸���o�9�tf���x�(8HL�S�Հ�8��6�E�U��8�G|���*�0��k������e��fPM�`N�R�\�