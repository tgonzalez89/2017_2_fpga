-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
zfPkzeDiuRL8srAqTfBMPVtdWKi6NklDf0G9/y42Z9Vsv668q9DRy+jfo8tmZLbYsAueCcc69Ngk
ywTUcuCXgcg1HV4SLT4bLwnNLsmt8AL/GggucZyCQ+HPWOlRYDHo2PiGUJdFE8YobGRrKsT8PHO6
mBYox+q+ITJY7CHHF0i8P/f0jS+mBFCEFDDY7yOR3hPzj/wa1HhtpVZBLX1EqyNeai5omiwPdAlt
1h5ZNeJjsSaXyT3EGApZ7B/9mlWP3U2z5hV5hwb5OJpyHCcxhzNpltyytw30SZQZ+h9WmaUV+oq/
UMh70YVgkItXGr4Y9i0OdzJWJ3QePdJyx3DIYQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8800)
`protect data_block
UEEvrTXE8UA68q/OmR+m87Rr78qQ0x4oUAz1IvUw5no1sYKU74ksHuIvUYWJoZ+1Wqk/uoNftM79
ahDjI2dygy09zyykq8Zn2vtSlpkg9ebeLT5zHmDTH1o1dhm/LV0ZbfjVeLRw3VeCHEUPAOzuL6ir
wYW5WC5h7VkZZZSR1gvOxVk9WQaPIxWvwvs0A26mYX02Qi8ieRe+GbzNVnr8ebZdupOP74CZTXZS
CUKbs42l2JfCoEtV4b6Kw+bwQWMgWaQXg3P3r38+JZlExEpgacuZMg5WZSTR8b+w9qkdMAfJqSff
q2hgBDTsm1o7Ir1GOFGsRuEfC77P4LK0f93g0Dx0MTwM9+4qpAXqspjRkwOIO9nactlS6e91pT0r
BhDTT/H0j071MCdigH8HeYF4eu0QwPiKgxw8RvURDSDLcFuX9+zfsIWvsfMtOUj6SvrfJ3VGOXzZ
3N3ePgj2HRos8ZyOpotMSExQmGp+0uUO2CMY03EojvHJ6Mx9mue0ENAoR/iOmmUXZ2Ouqau9HRMF
EAzspciPDyRl0CSb/IvkRbDTgMp/yEEo/Os7bAdy1oVmHCew88ty3StpLtt9TbcSn+ws529AtEQN
jkivDAo2moC00U6+9M7Js2GVJGE1/1qN/Pw3AirSPdfBDs+4KCr0hD9+8mnYm6aCCgT87leEQTDP
MCfMuuIRk5OWW7ZOFgHwPIacMSs0mvcaJb+HPvlBPuFzGoH0O3asbM3m8C1FNNj4vvp5rVf9dTj4
DZBfo3SWR1K/K2EqKpoiTACiGQElGuh1cJs8wWlg7jVAZo+dNfsE6jObG7CzsI5ibZwIue4WSU7A
8SFQhy30q5ZLVBRlEvop7MAt0eRWU+ifSkv1Tw91xhDm4FcjBYJeDIBew+nupFsiRW9hvKeUfiE2
FIagM4O3QlE8kBkzLYDqn8morBoPtrVWIpumuIEhzeaYTpOwuNemKqBNmm5d05lEz5pqEbb2wvIg
ZJm33YIRd6gE37twVNEBDKsmUL4oKXgEilIsnbBLTriq/3Pf3kZn6acf75sKibjYKWuheYvGXabu
F3uFWufVHKULK8Vr29IZJyCR/CK6TZpNS50ZfF/gc/xoshh5/JKpTgn3b4hNbrRgDMnMJ93S20e7
MNstmFRWQWE463vdfY9TQ0a9Zrd/gkFNmzrbv70Ig9cBXb70SmrxCAwmuo60k1LN0J6TJnJHqCik
FBpAhz/2VLEjEvCeAB2x8Rapv4IxvmlMeflHfKQ12P/Ddsm0SHoNKKfXnfZhn6X99gucpy8rhSlb
uiOeta3dUar0Gw3MqTQ2nHMKXBF7Sn12ggAIuOSVJBMQr2KXx8geCtdRpfywxSSC77NIQPfbC+V7
nnwsYIq9ObW/VUaa5Afros0vFFf2jvGSDLxXQjgA9fpOD2WwqzI9Kig3WJoJIJfoGcafikSx1Uyl
2LsVJvmyTZEYTC04IB+fO0W2W8ZNpLqUGyxMXXDuP7MY1mdvrGM2btKcmlQ3DXFyI8Sk9YIuPZmO
hCNPmqgIjv/nwcXu6GVeh/hgQlwCjwTMf0Zdvp/PVsCo/7eUD2tHqvnD5Hu3quO/r4/O7eT14+QT
d2Qdxf49AtuNVmnE9Qyec/7AIPYW+jpK4fxL+n9T3ogi+6KNqJ+h/oGwZ5LdDJavoUg7suv6345j
NnuPmKrm0EzU8vmBc0RysEmW9sZFswquHATjCRyZB01Ugf4ZGpF9X/Tk4W0J7ntXu5sZPp7WVP0l
uHE4Gw8/LVqOxC/JO+fb3sUYkibuo5KzhoihcfVfU3mE7TvsZpCBpHM3+JxJ0QP5Dkiv5glD6TLy
RKUDdFPmj1PwyYLKhMP+M3cHCYCHMrLnQQR9Fr9GyP2Eh5cS8Y6jUsuYgQCZn581KrETNr/Vc/++
W/CGVF2evz2Q9tsQN5BkOkJBsCN8J6M+uCgh/DjJgylz9nJUzXYLRNR6sDOQC+QwNepScr/X76lt
P/xqawbZwoOk2jZPWXRskXXjoiOZTBRXYb0jg6ppfvGkuhi7mxX6meT3XVWtOnd37JWcdcDgQM5H
/Yc13cMyYNofIvoLHGeBKeGMGGAM4s88dtMrMqxYv5Bmx52opr6uUQAT7uFfaqj5UKSZlZ77PNF2
k9etXD2a/EbIZaiXwKaFafIOXcNZ0sR/ezKfGrEq9LJqTBd2Jg/FXShmLGtNUX3UE6zNJI3y5a1X
DA7mAYCSk9aDx8Ok2IRvEQVXs3n+dYy2PVZ82zyG9MgGLuY324T+iu1HlVlG9rDG3TTfWiEsX/bi
bSTxVIWFekwHCNSsJUEUnX8bvVuvMIjlKLcx3LtHJawYdHKxsuuJiR5QxMd4iGeUMgyZyX2lb+3G
0Ue1BPdXzOuL5WkbOsnUSurtB4RB5fimXI45Vbd3l7IPKPZrJJe2RlScxuGuGh0/lkFfus+RUSyf
BLiIYHWrLekikXeC9tKT4GfzsC3YpTJEY0TTpcSm2uRsHeAnBrZs9ZOVwDN3V2S2dkiTUI4s5QUV
vl4gFwkxQiwctC71H+66Mrdgrdz8Cv/ZtYJeqePLsUlPZ5ds70E/UZXIuPRenOEiEhC86chohwiI
vZfJrp4xROQtjz2tAZ1DvlMuNf67im4VXCmFSXqJJHVMdA0iytsi7Lj9e6PKRapfh4dc0f/6/SLS
GT3BM2rLLqOddUsm8DDigu+ZKI2p1ydK4qQv/vL9gpcuUqSx6uxqs8mbv7le+KqiAJqBIbWZrbYU
FRM1e5c9SwG9FRAthRum5IZO/VJXcZ/tAVzg3pdHQdIIAV/mslgcen7GxZLLWGZWJXAJMVT4jgzh
z0L0CqNcj69ew9dQ2DLuLEGHXqYANR1DgcPIUAMWIy7YpHkh5vy1gQ/JdTOvTav6vNaK1TBK1NtZ
Z/OUPsL93afTDNRti34t/c2IjxZtu17A0pAWBzvFUCgMiTRe7eNzcMzrQKItDfXDQ21GXYrjZU47
A6UOJfNcAHb/mWLJuxVCd/zoZhp2PwKNnCUFeMpeEqHGn1Vt7AmTOOyMifGJ1JPFIXnaiwdaUw47
HDQpLGCMFNzFkOzG4KzLbZo/btRscUl0RAH4aKOo5p3CNSH1FZohEfuchkluIGAqPQhD8wYQLwi4
6ocWUAoAUmpIw0+0TqFDAPB3dn3Q17kqxNyJRwWEboIkkbAPnomtz+b8SoomP8Ycl4kDcJ53sNIJ
yM3w5UYAp67L/vtKL9kkN5zcMa7pAiP2nmruSC2tKvhgMalXrXHGOG0Gfv4d3+S8vaDqfWCzahqO
p9uts1ndGjmsdvksCKI5I6uwaG30yPq8tZeKesNiVSiIOuEiZIVKP8fNa1NvKpLLuU2q0tbcv3tq
0EojFim0WtX8omQxwRMwjUmU2+aqg7zzl3+tTgowgR86kbL5Vi0DO5DAChRXZNirHp+0ZUO7tv77
yOUiBAsLzttwVMQvbWnY8vt9pszOt6VM1qNujjWlSjheoaAqLBthLv1PXQHxVwLxaSbxf2/Z07qh
OpSYJC7tz8ab4lBhZyfrfrIIifVNb/WvE0pAfwe8ugQRdHWUFIR1qVT6v8u1xEYjCTidqu1JjT4V
jXSgRn1IP7mtDib1+tFYd4GQ+NwyeX7PytNbJosj0Ug+nLNo2LiDfqbRriT+fe8U5unsnuhrxRVJ
o1iejzmj83V2gfDeKxtaAJp14S6dbYyH17igp+7UdxWVJgAHDrCqU9bL5xxJ74dsr2bRY7jcoXQE
5oBi5x7CwXO1chdHwR/aK/VJD78jOcTotSD1Kdzct3Sh2t7edJ0m2pB0FJvGCKOfKmqRdkg/GwxB
tFeE6JxVs+34z8WYmB2N+byUUp6MUBLsmIWK6Bclea867KyrAAWH5yM8FPABZEXUkzoVprTsqZJ2
HnHmuaKDEiPnxsO1XkK0YjIGTB208LX115m7n/dshtOq7FMsfveV4dXM0ljmcvxmMoj26Jg/f0G6
RtyIeOg63pXKF2ajm1hmS+sUIgUX4RMmbwxTz7zoT/l0NFmHjgCA8tV1GaTR4kE91RWEB8xjayel
xJILx25PfKFrY5lidIkiyjNqXcZNGH77iaFMCI2QOmikBTOxzxJCs0MZhZxLQERkpHloqjBpWVwA
m5NJCTutwJ1RLS92mjrIieDeXg/S1sldpcjfOn737KxdtJFfjIDbCSWNlFCawQj+njBuaXLL0iZx
+xR7QyJikFVNueeusLEMZAspfl8fbYY3i6bHzUHw+/srRPh3+oailc8zyeTuUQ2OFDACHsBZwG8F
Xu/Vrwj657Y1b0AzivZ6Qq7xixJaG0qSVwbylO3q6bXkFDSSSn9/jctjTxldkn9U8l64jbWVUxBd
fBifzHAablVVxh6C0gYugajOdUV1rniQNN2wDBsKj7X61Y8KiCy5fhfwtfrVL/fpORVW4/j2SgIw
+y01MNLGNECyMLLI3+C9nGnDZi9LmpEf+2j3Xd//BdJOvsu2AozC5pjXenXOiLAUxOIlOGx48uYv
aoEnkUqxs40FI15iQB2ke+FHmuSqGlMn6ek6ftcFUuJn9br/RMH2H84bNb3G+zzp2OFen/efL8xI
svQ+MbqfTDUq69XD5QuM3W0rK3aCTWPOcGMGOnQxxVe/7XwA8JQA2kSmXg7PQSPh+Hr/0T6jrZjB
cHT/4EWdev+JgpII1OalBdfxO6BI+fhx/IIqsbzXHO9svouuFVaToTRf62jxaJU2nIsFgQgcIsNP
IzwYN/MeIL18vuTq2au9p5j+KlpwdwMyf8yO5eqqNPCVcgCakhEvvv5ipGuvhb/zkdQ+xTPM52HN
YH+hc6nUF1BqkDIytjQOK0waY3Pod3CmJycTg+8cvdIkbo5rQw/U/WgtmPumhfV59DxCKaeyoP9a
iWvOpyV7TCMUhBni3dIAceTI5TynX7xbGSTho15Xoz3FxZBGsFPJs9BLJm+LEgqpJwUdgVU++VYv
D6nwL+ooyt3rTij4KrrgAODzrhBhKCyIydwsmGC2HeG7Z68N57UoGswJXomlOJYwttA+L2fKFPUj
e7hcgyiPrWAOeCj3Y5yzePH0F4sUvlr9b+gfwWcvMTfC9kZFNvBcOV6YIwxwW4SUQ/UEHnTQvV1A
ucOQ7vS0fU2Y/8Ym45azQeO8BakOwp3J4V92X1jbSHfLv1UvM4iHXvwxDtWaeToxXyvcMkFR8lyb
TJ7+TsasRfOeT9KBXIpXrfaJrmaRlM4MeApe0WleivQI28+aFljTE9jmLpGUX/YJbEdVWZ7P+7xQ
eaJg7JLRyCvJddz8wSfgchs4XiqdxWFZGK0AADuH6aqcd2+MBHZYAZ51ZrJxWLXNdz4A1/fTcFvV
z0aWWOhYwbqn1NdYeKnuF16nOay3RRonYX5diz+lLhRQ2q5/OQJYdszjRdIIGCahAALceABk8j2L
n9gOPuXC0osfAeHd42INi1TU1X34jC7BNme2cwsx/1hCqcTLuRo+uH7V6nKfAVNiAyySCZOcd6ob
YNAj83VTMFAVBcHDkEVABY5KnWVTqbtDQWdFD+YQsoiZyQ5q22unjCrRYUNXUQHd/HN4vp2i4XEb
S65YZEVcDpYn1Zust9+5LJeeYwFDrT0WSxMbfQURZdf4vH1AfMzVrY+2JcHgG85UNB3WCfYMCdEV
YusFxOgkR2RySMxZRzNxMFGo3XUlgNWKO7WO7m9uXJPFVKmtUmaJnzSZhLY+9fZHSSoxrGKsWutN
Em5AP94LW8OV8VAH4Jxwtc/zZWlAA4zmV3i2GeOWAJ3fqsqgbK5yaSHVuJI05kKxnDobtpJ2T/R7
7n/lPMMnyd+QXvk3bQaxDp8Jln/TkFmsKUEcgr4H84XcepBtKbApMxW1MUeUJsq4DuW+9IEs44Y7
oJjLe5LF7tKeGcx3NY+OFuSGNcobNa1YUwzV8KdEBha1usx9tGOnHm0+Xd0c+ZQK9JWykkeHpG8f
63/k8YBZW+qkPH4zCcJdqVADoH3vGHJmpRMSkVZADvqo/EcUpmVLthbAnSCtYzg5cfs+DUtXPL1b
C0C67CIgvN7YHo3agdr5ten34tczKhTySKC2Ia01trrJrRWncqv4Ol7xPO2P5hkekgFqmSSelkqv
EoRamGWJO1IEr2NHLX3GzP2RB+OUKG5/tUpV9XOMVjfYCf2IM7xL9HcqFcRQGgxUvjP/H3/oMy8J
MmYlNUDrwELwTu0Ywgwz+apBomLFcIswzjZZXS8h2xZRZCz0FD3/BKrGJijo/L+nCEbtk4rRkDJ5
mwdV3V8eTiaKj65AR0s4H0KWHRYUPTr3SHyh9vdPtm0dkuDKwtcfceYv8eULUrEtGXUr52BE/K4y
w/DJmY4bSYLKMQEZidw8OB8hfD4Z26t4gv90d46e3K9MJOWBxuv374ecGvfeeISWGsUNtwjyRXe3
GQbMy5kLeYiqr52nJKC6jOVOIgvyw+LKUmiFVl0NSx4fDdyozACwglvA6ks3KGJjhHM72l0XgZ+d
bFn7n8snjijwevdkab3TMMB+D0dgNJCD2wQq+kYKXqG+cMYdK/c5HIvOZUFJHF0+qpeWdbA6fjCF
KcccEaB0Kd6SVeZy2+3UeeQK4315ogqX2zisTZqjtgsHoDl858ylddIXovO3jKlIRnrMyWB9HKTj
Q5RAJuO4uw2BCMBH2eXkokrO1JFfSwRwAtSxdrOIgtWRgDK7/SapJ5UPfwlmoV1il2239/Kt8/7e
u+KHoxygKcMfRRbfEbpWrtx/sLo7RnT9jvfFuBr6RGx/q0P1DpiKQUFfzd4Fa+8Xh3W6ABG0WfwM
VUYgTlgeG1J42LbnqfSZf2LxD7gpXD3DY24VHC8om0tMvvDOdt49bRtypcPCGMHLcGjrBzHQFTbO
VXSXFyIg3/3pN58uFxudPgjqKsNHbJ2PmmH6NCyOha2LWpzdDXrYydxkc09BRoTv0g6tmpIFueau
fi4Olssb3MH6EJt9wj12NZrdfpSMK7+lvE7Xm2pIm0/ceIIIn5NA5s/k/KXdIQuNX5UZY1Zn4Zvw
BhTQiKP4hYmrohTSNPII6hCekJZ86/yQBI7IinOnbPOzJ+uD/XTCmpRR9JpjMDtFi+DrZjJTKuXr
UdW8re5r/4EK+yRKFhbeNYLCLvKoWS5GabO9MU70TYRYSFWCy3jrt1dUevdPXN9JkGpIxYwMwOtW
20eLwptIgjfy09CJ69m8UK754XdOvjsMr20ITXfKJmV+DdleTSNkYpUZUMAtB4wqez/xd4lgkwJX
ELPZAnZx7VWUg5th/HSm49Y1HIdvMvZDYODqyy6iG6AqkHeF+SOJAtbYvmrXpHgCvZM44fhrJddN
/Yv81M1G8t1UiM6mVXHLEsljm+3ab0NO6W9ixwHW2Uw7FYDbm/rItXp2ZabMFQTRNCX7pQnEerco
IteV4PT4KkUga6ABqjavB9iZ6KyhezXQVocQik5CN/q2Zh+gl1rqmV5scwTJBgqjuBH3PX8J7kmE
/CFlp/Zzhx6XCZ5Z3c6/cRM/CR8UrRfwC290sq4B0B3GITt1YhiWgziT9aQZw6Sfe+SBifJTGTUC
40Ujj8fLRXrkx3LQiHJM5NfZS6uYRHDfh7cghySC5OTwGjLWleq/DmHvk9ApQpZJ8vDODwIrIKas
AoB+wV0cG2ZNOI9PlUTa/3BSRphfJeiehNQ3XXTNlGf8bnSeXh6kQ/mi5sY3rFfafVrE5gX3xd/Z
h6c7ioTEt8tgEPzpgwDi4Lp6aH7XL50YK0aXfZLJ9T/jmKA9Wba3Lqbk/c24bRSO0RMcDPTC9Sds
TOKjLbRtSx2jFLEsz//Xhdwrs7NsW8JlQcuBpDluu6mYYQKHRxy31HrgUg9OAzvHY5lt+E5REOM5
ddtVzdB6TgoUzu6qkWsKrlMB6+DomvnXwl/LbX4VB0tA8GVt3iSwDaCPywrgxH9KnQWkT95uzPwT
usmdcfBOX8IMGSOZ+HKJaQdO3iocL5j/Znc3TTgxduJPBggdKv0ZxOXec9BdCv1/hR0IiM0IizTT
FBlULe32duqEGMasqln1hCCkqb6iSqerO4vLKJTrEMY0IcJ7pO8IUA+HdUj9tXU1eNTSNwFQSL9p
lbJnO0mF+TpPuLusb4su+9IxyDeiqV87gbqTEzQSVevNVs01KvTrif1+EeI1AvEOlqoadENIzhpF
ygtvAvDL4OZJZUvHC+Lj2bDdEX04JJZNpjNLtghZTk6iTTMjRZuc3owPMgEclkoHPyLEmqSwYHdM
njr4MMnKCAVvK+JKL5kP8/j1e+9lbrBEfsj9UQTh72RQAT+xjmt4DkJnVPZctNH5CcDAwxEwKqqf
9yGSgObm6h1/tk4SeysjGB1WxiNvqC2WWAlu3npb9QOZ6s7MySfvpYEy9Ona0n8JOKXtTXDBuUps
i7wXPFY9trWqyysmffMhdWAJ4iIGt/4IapQaTAw1nB1biJf4PmhGQfcN3F4pm09e7KMKguNaWxBu
vfm4Eif9vd973P8IhAR9z8lTcpOp1592TXEpFwPztd3luYVJdmSzdLsJCVjXxQWO9bj3+EOp20ee
Mnm4wTA+eS7cejSBUtE27UQkdNbzKIGkU4z6nhFWf9AdH0aCuCEuOOtkdorbLQPnx0sBTEwtpk5X
Ic885W9dbWuiLq2lJE6JN/seKLnJAfBWTX/GsJzP9C+QZLCnSYN8dcoSLQlk/zDadA5ZqidQVrLi
W2QNpjOgnaqo1TVL/rehFdLRIxv+R52vN5Cu61MdPSUzoWQhErZTGNQk4IWBaTEmScUIIaqkQse0
scfFQ+DDLF2HhwqlnqR1JK0xMaqj7VCzTA0x3b1Sxsr/0aTMMvfjrB0j8sLnJUf/5UNM3UUsjcbR
oPjDbAT+/ezM2wg1tpFctl+PaKLFksm/UzL04mPSTc4F+wcOt6bh19Qdfqg+NIqsqvpO13c/uIzj
n9ahrmGThM/iR6vTl31ri1Uo74NXgAKRMcHzCyaf7gxq2dGlnX+XpEiQIeoajlygH3C8GL33uin+
tVHcRR4Ghrsv+aBe39TO1a4voKJ2BcZUIjH3mZgA1I2vozkYT8wp8TOZZjY4BwoM+l6ibTStom13
X255oM4ymmIcQ3QorD/r7VksUws5HACS1GUDe97Kdag4ddgipvSEAWGcdmMnIRo/YhkscpWIc4Il
PZDgQCuRc8AcY2up5NsRapKy3OxOTv6u8u6kt9FUvkthGzNGUzdFWlxJoA7C+olhtBrZLNSqYK/l
ptZouuRrC9goEa46/EnY3a6d6eSBL03tkSgQlrTpnxKtvlbDgkM4AEkS62S2H0Z47BzJOkJoTM9U
JODwsVkqdzcwX9tb3wul8QJ9/CJl6xMo4cdvMDhh0tXIBAVyWMQeXL+H8c26t0jsog5QJPRo8GmZ
fpNNbZx9iNaI8xvAKuSE2P/WClkuFK8wRRYN2MZG3PtJ1PuvsMAyHa9+3QUAkXz3uaEmNhE/o7+W
tJQ3rqjfspaYJpleGOMLlcnpEcFWGs/1iDScM0JHX28fQeDh6m8gyxszbPL7qn4xNO2GnJ8kOp2k
YP8Ch2B1RpPAgATywFCJOL4Vjrv85eBXNGP+7ry9ar9L0lpLC4DrcQx7ulgE2psJPwqjxwkE8Ukn
w1YiP+riszk8jP4fRav6NHLN7p1U+HrvjubUuHTq0Gkght+xFYeXYofK/yzUc4Jnh0HpsKje2DyW
MVJm1pSs1NLQsLjU39wIdguLf5yBXhkQKrnxs3MliRIQjDh8lV9XRWJ9QN+38/E5TqMDt3QXHW+R
Rs0X1V3Wk9YXA35P5s7dotD87rGteuspdUyq+KxrgGtt96EIk62uNf0HeHaYfBNBW0ZWq6iGRe45
16fnryMrW0Z+BGmASGxArU0TCguqTgSuJ81w+VVKkRLqJiBKLQnrsb+0DbSieoAC4wE93mBf0A6H
3WDVMAigUXLhDfMmKIE7zu8oswH1fGnoaPKpoclmUuvvUaw5K8j0rb+rFULMvCGMFdPi52wA7MOT
wqz22YjsFvvDFoCrN+Pb1O6B3Er3cEt4AdOsYwvNJVkbFNveyP9oijo2wpI1VD/sVHAOoe49qSmU
thB5njkki8jvQ9UFi1sVufuTXufUVZp+KuIlUIXR8Y0gLsZO4V3vixguFqB0ltjwOSTFXq9ppCEZ
UQXuBlXc4FFlyuBUyKEa1ZVpzmaMZD3QwacD0XvE36BghIF3zvxq5X8RGpxib2htVLUw0JHtuj4a
Xj1S0FDQ2ILlmQ+3G/iqAlBzGGMyZ8NPs2VqSnPp62ftYvaCWA00tkrQ9/+qTld+7ubV6Rf4s9p7
lp4XPui4tcGLzikt/T4Q2jhSUrUaXYthvm4bF3TkRTCczuEj8bRLqj3SrDTSyRHpDvvxouuIWHDL
ung+mCBsJ4U9E9ELpC94yG0ZEfpdkWyuE6FdYHWIH9hytwrJHIm3TAbVb39NBiLUxuaWAswCGuD1
IldKgYMk9lIUCFEQzamKeo6+AT9frRTm+z4iVmH4Oy6yOSkcQrgqZo7VltwvwFj+EMmyTegQxydZ
2kYGrHc1fiv+PjWZshvNAD7uQjQYGBc+YMmyqlK72VTvqGdXK63AWTD7JoiwUBCeD7acnGQdL1Ud
fpRZgwv4fWzxyIUysWy66JPMem4TdB3rr+kYND0L75SwtiP5JenDI5u6FFNJOWm7zQU1wDWnCPr+
peoYXfoIFwGfLMS8ZeSynea6YNdKQlUX9WKM+vDPrHdHVxd969SSTxBHRYgQj4UZqje2QGOBu5MX
uuPqwjE2sfhfi+T5zNTudBopDVq4dKLh41KQ5tEtUuEW9si9pkXOo4wvI4V5/8SmZNSBrR1URoZV
kty9wRToEWxhh2Uq29PPo7mevLZAtl5fehOu/oZ3HRb8+BqSkXrztResqRmUJN275Y1Nf7YLJR9/
iFh244RENTpkQeGRiBLtXTOw2e63PF2HmiuanPCNSMMcskJQTdZ8EmILnKdj9iOymjvSDVmq/NTE
VXolKQbAg/NMtti23Hxj3XPRe5wDyvH1b0tHm2fvrk2GK5hmcBBI9Guqzk9zzkn5sb9BmHYjLuJg
NYKzAMTU2jAtCyGOkQG7ZTKOdGYeIDo+AmxAvLn90d9Bd5mJ+t2H8cvK1kfL0hyVzG5EgFX5W/C+
dI5EDjGbZcO7Vj4FU95vvzqeSf8FvYtnv3gA5Sd1cgDiUbGMOhdMh4xrVfbjAx2icxf1VHXUZZfm
gTuGZ4U3fMjSy3xk5bJhLkIkunR3o0yuzRGe33paCwz+EmsfbQRpC+Ix1Pg4xmX0KPH6kEYlNqOT
d6JxhreYTG3KnEQ09v+s67F0++/yCvTgVvu4G4eeXaDMg4bhH2jLL50wLvScxt1YBNpgvqh7X4C/
pv5FBsEwgfYDiV0Mrb4z4qO14dGfRstQ07C66CGzU5TQFW9+sNalXzc0I+3R++VVUw/4UYHFS7cu
vxlTZDqHoq5FplmYpEhuZjAgIEwCLSrYTnf1NBjKbw+90JI6SeIbdDc022LpUhG3cihTKdKms2Lb
f7fKl8eck73uF1qICpC7ljjs2SzZzott4He7ALoS6Fni1w6rgCfnlNrFjFeR1xmCSRjCOJCM6t7+
vnqtpav9v+nsNLg9ZWQKlAQ3LndUEN7nnDT52r0vbj09R5ArVkdtv0GK214AJSIXZyTNhmzNB6+Y
eqPZ5A0vqDovk6hXqdXSm0VlnKicdW06+Zzb4OQ69Cnvj2/z2TadfORq92ntfrBuczCro21LPUQZ
PEwpS4+qiV8AWsg2kKq0JTx+dWuQtw==
`protect end_protected
