`timescale 1ns/100ps

module tb_proyecto2 ();

	reg Mclk;
	reg nReset;
	reg Data_Available;
	reg [7:0] BUS_IN;
	reg Read_RQ;
	reg SPI_MISO;
	reg [7:0] Address;
	reg rst_clk;
	
	wire [120:0] BUS_OUT;
	wire SPI_clk;
	wire SPI_CS;
	wire SPI_MOSI;
	
	proyecto2 U0 (.Mclk(Mclk),.nReset(nReset),.Data_Available(Data_Available),.BUS_IN(BUS_IN),.Read_RQ(Read_RQ),.BUS_OUT(BUS_OUT),.SPI_clk(SPI_clk),.SPI_CS(SPI_CS),.SPI_MOSI(SPI_MOSI),.SPI_MISO(SPI_MISO),.Address(Address),.rst_clk(rst_clk));
	initial begin
		Mclk=0;
		nReset = 1;
		Data_Available = 1;
		BUS_IN = 8'h00;
		Read_RQ = 0;
		SPI_MISO = 0;
		Address = 8'h0;	
		rst_clk=1;
	end
	
	always begin
		#10 Mclk = ~Mclk;
	end
	
	initial begin		
		#100 rst_clk=0;
		#10000000 nReset = 0; Data_Available = 1; BUS_IN = 8'h3f;
		#5120 Data_Available = 0;
		#5120 Data_Available = 1;

		#100 Data_Available = 1; BUS_IN = 8'ha0;
		#5120 Data_Available = 0;
		#5120 Data_Available = 1;

		#100 Data_Available = 1; BUS_IN = 8'hbc;
		#5120 Data_Available = 0;
		#5120 Data_Available = 1;

		#100 Data_Available = 1; BUS_IN = 8'hfa;
		#5120 Data_Available = 0;
		#5120 Data_Available = 1;	
		
		
		#100 Data_Available = 1; BUS_IN = 8'hdf;
		#5120 Data_Available = 0;
		#5120 Data_Available = 1;	

		#100 Data_Available = 1; BUS_IN = 8'he3;
		#5120 Data_Available = 0;
		#5120 Data_Available = 1;	

		#100 Data_Available = 1; BUS_IN = 8'h41;
		#5120 Data_Available = 0;
		#5120 Data_Available = 1;	

		#100 Data_Available = 1; BUS_IN = 8'h00;
		#5120 Data_Available = 0;
		#5120 Data_Available = 1;	

		#100 Data_Available = 1; BUS_IN = 8'h21;
		#5120 Data_Available = 0;
		#5120 Data_Available = 1;	

		#100 Data_Available = 1; BUS_IN = 8'hbb;
		#5120 Data_Available = 0;
		#5120 Data_Available = 1;	

		#100 Data_Available = 1; BUS_IN = 8'hc9;
		#5120 Data_Available = 0;
		#5120 Data_Available = 1;	

		#100 Data_Available = 1; BUS_IN = 8'hfa;
		#5120 Data_Available = 0;
		#5120 Data_Available = 1;	

		#100 Data_Available = 1; BUS_IN = 8'he2;
		#5120 Data_Available = 0;
		#5120 Data_Available = 1;	

		#100 Data_Available = 1; BUS_IN = 8'h5a;
		#5120 Data_Available = 0;
		#5120 Data_Available = 1;	

		#100 Data_Available = 1; BUS_IN = 8'h1f;
		#5120 Data_Available = 0;
		#5120 Data_Available = 1;	
		
		
		#10000000;
		#10000000;
		#10000000;
		#10000000;
		#10000000;
		#10000000;
		#10000000;
		#10000000;
		#10000000;
		#10000000;
		#10000000;

		$finish;
	end
	
endmodule
