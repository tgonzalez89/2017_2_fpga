-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Cymyina+xx+7Sc9ku3jQEDSbc8vdcfvbqrRyK6LOlAQK5sUkm3ca2mJxH/RdbbDm9G/bnAL3WzgT
OMqBeBCgVaEQ/B6gYrvR+EpVjCTcI219LwsD759BRwy4+l6q5t63rzhtsIlnX26As6zvZKczDHaF
jFkjjrkyJR8G/PP9dDqp0YE2UAcXtgMtIoKJ4ND5g3YoFGxLUu504GHNDOvU7mDG0C0PeVl9U9L0
ustLxn2xO7dp9FVS2uc20C7ib4uAG5hZ8RDDIIiUp83FVuXZbPs4654jqIfE1ErNRr0aMpvEobRf
jzxk12JQj2vv3lp0AFce7afczTu/AMGveLHH1A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 28112)
`protect data_block
JqD9XCnqfPFjtEWTrzZzzumXmz66JikYrC2jGyioswtGk4VOdnnxNyT44EHSRggvowftSLuIdwz9
3DdVbWHqt+4q7nlwerHQuEQf0PoXGpYknymqVD1ehcbO3sV876FCj7RxKye56ARcOGFP1PcTxTdk
BnOo+Pi2f798hqfTA9zcH2av33fXNGwoeruPtxlRuGuN99wDbktAALapgAACFr7VAjlTBVnUc98P
gt2XaWxDMPUcJ3in0D7IOLt89hF7Yza1jdnH3mWrjICeYOLyX5Im5f+l/jFW8oS27SzrjyeNMawT
oXhSkk6Rsloj/O4GIlOWCOtb5vNygOkRgmJuhNxTstBrGza/jmg56M2bWFcCOwUXUNEItOswrj6+
YnTEcafWqmCgQR7qqBXooUWyslt7CFHfuoTGDalvpTmJnF1pFb46umyickFQJHJ5fPlhG7NiBCJB
yW7PeM3H2FoKz63CThcPtGs0JN6RMddkX7h17SCOcKlcdEnTu2UESVGPJFOSJ/RZoswLnHBe8mlU
EnePA/z9wQeqvdDOOh7BZW/OhNcI3S/PVEVfZa6Ak/YyBMBzLtEKRo0OjkvL8QFsMDvXgaVWVykb
wr9X04Ni2FSFCRvLaHAzxj+gJESx/jRLFVA5XS+GZK4Ms9y1m5cWP3W6YVuL6YzYzH3m0BQOpwXM
4jTBDB0AXK1cunk9KoCjKFIjtRqZEpWvWUcuc2Yso9AkHkdcCc89xFEoV1GlAr5UFVL82xcZifte
bK6wEwiGiFoecj08iFYIYn956Q4D4Za9vEZishgYIxtJD6ifUc9Fez01YCSWUgjRnLBU4Q3TchmK
tJbcKgGZX6S+Yk/yieyiq7xKxX9ymLoVYbcMOmcHQmfSZOgIXhfLyc9H34tOXj+vx5JuJWtWyrKX
uLFHndvN5wBV7Tci46f/+hFQrhux/Bkzb2TqGDaxYodxRQE2Us0tdWHxFd2OftUsOww/tViXMQnH
sJJ+i0t2wSxmsgiPgE22v7aiVRHACwVSjGdNSv9aidmzPEfiBmk5g/MJ74LcQFg7eVpDONTF7SdR
4197/+aUjMSYwGxej0MMGTk/bxfQYGJ+LgbdJN6ewmVMzOD+m0Pk4XrtH96AT9gh6hdh+HwkRA2y
2oGP5kKzz5DjdEewv1uV0iYxp+9o3wY4To+8bedbhPHgSZrq7C6vCG0d5eOLyuKHq+tYeDbpjM6u
mrsShAZBgA3rspvf3n4+rbQgKPqVJOqOR5lkEjWHn+m4vB3uW583xQxk5/v/OXygd+INROXcH1nd
B1wpEkVtHCbRP4wOlTLbG+QIn49wgmt0/irpP9zZsuUNVR3HppwbVETqaPZTQkkkx4R3h/tnvfd5
nFigWzHnzTS6fVce0hbXNzhzHHFYSQS9DeXcEoYj/FKiFRaG2qUSSy+mm/3zNBAaqsyQyjWeeah6
o9852YzPW9gem3h6WaTj8F7O5n/GcZR9zT0+g9tmGTsBtNmKyO2UWlnmKxakG+yb/7WrvQywX94O
ugmMn/Ho/DCLe/5kkDTYO3us59aGT79qo8k+bXuGIPIjkk0KRaaaK18+Gk5awf+SElXZYs+cBpjo
0jcj8aXV1UbKiJfHNMe/jINFN+OAV8rtNV/Jla6IDICbSyN9e8OFWJuFD30M6397LzI+lemO952Z
KtOD9+jLWB3FItbzAHrrwgol6Zk2KDQiQWHeIlPEe8DerCc0ffUAe+5YrTAyevA1J6QB+HnLFlzw
55jwCneZd9pNDuXtZDe09J23vpYCWgLBAFjAMCpmXtpAEOOjCGeFR/xjn63pHQEyMjVsKXux3EGv
FCUG3IHP5ksjBuKRAKepTgYrZp/puxH2Lsm0LfK0/iqtkqTCatHuLoQgSA2wXIOdgk52x8k0YlVT
sj0Rr2YvxLRRXq+Lrf2diXLP+XqYqhQoV2I0wK15ChnPJs/k8Kjm1klhC3ws/obVjYsuiUlR9r/6
gkCJUICrFd/bKT1SSRmscN9LFc7S9SThvhFux/c9Z6lnqc2w+Ww1WrNmtV4ZoEljRLqe3UZIJjwt
U0EtavI66Rr4D+7TmgYecBKv8ctanTwd4gN8mXYXJWyBMyA5jdo7mArVHa6tl/lSBN15x7oHqNtT
qpz5RtDgyfJEI2U6dXLpPmnHKRHx6lQYTlirdQL7+kBVDbKu8N6yXuYb0TnAoMVnFqEWwyebT5iL
fo8DYqTKpb7xz2A4LfuRbKvtB6835FVhFonrJChKlwD6xdXJw366ywGDNDhvJrqTFeCN1kE6T0Pl
K7RB/OUrZ15EBY1aY4natwAa/soRHGFTjlyynHU2PWRuEl20Mx2JT1qfQua9ftLzUaYJiqC9DH6K
ZB92ov3ypd4e/3fT56noHpFgc5U6Op6rySVdOo23ICsymVnXttSQzAnrw4tc86gsnsuEWGe5LhxZ
o5HeUlvwogRMkOSO31TjLQYToi2Mvk7EZ64xvDlQ7uTbyFHjeyNXW+69bJ914T6pXx42w8GL/Ih2
FNk+pSw91l7+3BzGKz0r9ifEZD/cTjpmlj5Qr+ypYO+OmFroezYqrjZ6/y7V+s6Axi9l7/5XbVh8
mF4sqho0u4oTRHm+XYIKJKd0L+XwOb9B4BjuFETUGjZGKd1klCIriatrW6QHTC+cAp2yw4lf86A7
uzkQZeHcEsPpNq88LVP0WwqDlnx2LDuyJ6fx1+XsfkLVdcyUdhKQ0fVdDW4XSUQR2mEfKEJ35A59
+dHHLxI+dDSK6lqvLWHfrW0cO/7/FnW1fmG84Z/f3a9bT6weWJ0r/+55gISfrhm4X5GkEWpCpjCx
a/uHANRjy+dzwVZjexBke4S6qH43hlzQ3VYFpHi1zNXPB0s6zdg5jeczszat61ZX/87pq+KfkJs1
0dAqJ+m8rzb7UbTdkhIkw99Lsp9/buJZitvqB5oCJKpbauJwnq+AU8eBGXySpo0qewawrNUaBiq5
NyDpozceufxdoMXbSnx5MLqqbVJ5edC3lyotttbzA7nBQRuHKSqS96PzorkJWAOB8q4bsX8H/QdN
yKYSLWXNTMfHgzJ/jfQo4Fu1rn+6xLObdep5qOh/+z7yy59Kb3hGgaM2ckkqJr9hVEVXwAm+kGJN
oEuZVBL68qR/fCriHEMCJyifKOT30TjIy2MbR0OLG2g82xT0eh2s72pE/3z9kMJUsIyz++UKqEZI
maqc1HyF9NMxPDwTArUaByhM37kMEl0wdw0Un83ROhDU7eyOsaLUUAnRZj92GuSCuZgZzzOIpVIm
7fgRXvFHNMYg96jLpcGOCkX8uz9eedDc6UBZD7INfckzt/YT7Iu1DPosHKCxa9GNCjtqGa/SLw4h
oT8BJIHnMwtv0vZ1M6hC4kKvOTg6+FeBQx1I3Vp0MBhDok6E1la7cgvcbVxcn2/mfJNT/k2DXX8d
BLq9vGfIWv+m51b/YE1SO4PCGGlUUcWF+gfbjalahPy1lcQTV+quHKMVZPwSZo7y0oTGDq1+H6Ue
RDORh2lJ300F+Xz02aSAU7lgUp73T6C9Fmf3bovdUEepZmMvdm9DsLYBrfvAXg/SRNBX85+KO7Xy
DcF87+0AOMZQI/dMxum8klsV2XswkVtVaWwGITFt4JxCq+wSgMnaoRaHNX8xZ7ktv1UFTgNapJ7R
xrwTSsGRiDIkSoTyP9v7DIskRVKo63jWCBnZ2sxcG9XX4fxuZ3wmo7vGy+ztJcgntwIgBB17zgc1
91zgKf1w3G5XMdvTPKHCIGlcaNy5b5JHH/hDHZ6Xhs2iTaqCF75j8qt32TGARDVKXPrmMDQi9kgh
M+Ckh5Y3nFKDxJWlIoSdlHoP/ZsJ8P1JMriR2S6qoSW5J6/Gb0R8eY/nPidFmyYPfbmJl4CwH1DH
ELfI1N7KqN/6BfQXCn7h1oWaO4G+qMTFNrIl87mm435oW2zwniNZsJSfHqkXsKHfLr52fGpQhYWI
ua8ZwR+0mRq6OjC3GOt6SHBk60rlIQsggBPIImm3mnNPPzILmDWiqVODgEFjiDDF5Ey0hHIzyDU2
ACsRyYe2V2j9FrOeFykbjw2HGzZr/+5O30cvzDoH8J3jLx+70Cgs58UB2fJFo26em3qAJkpbwv9C
ZqDpyObULntk8MhbDPXicm8v2DVt4fnSFnQnR0smA/16FfGI1lbKmyDKgSq61yJXhYdVFZ8vWCwa
tCyW0nR2OCLPftqMJHvX82L+BQn9XxM1tX/Sk8Kb98U/80E3lWeuqmAuPN9ezXA50oB9vElVhcNO
NARDfPD0e607lvULD1MvomYF2aVpEsNbg8H791f3IOpb7fXxWbWp/WV4xKzA0a6NckKAyvLkjal5
HgI8BeJwXReNio4tPW5/dms5uNLWzq22RpKinPw11tm/sG+VNWuaFDFuByh1TtWizTlLGYifDQU7
C1H154LLaHl79TG3kpwvNWyqvdZWF7j3Kw1bTR5O5bX2uJ6ZOi0T+5hFTOOs2APPpNXGxabZTzYH
M7vdz5UFuZ5W2vOsW/olhIXnydUZBjYy+wNl8GsUNYgrag6fLUAljdu8raPHdiGwEr6LvyjaKRM0
P3UdTnHnQZUZ8v6KWi/CvodoVleorWmt+vlXku1M5a+9SrhZjMyunztQA55R2T1RKsn6Pb0OeFZ6
78i/IydB40OocF6ER0JMj1I7B3dUFg573IU1jitYrPN/yX86NechR7g2c9F7EJ7170Ukq/NRMCH4
f2igCt+IwcMm4KF0eKswBYgW0gropyOZuUQq9tlkmqSWh087orMwYqUPnDv5xd9nSdk9+i3L8vOE
Gk5DT9CpvN+pOYWn1vqdFHEQr3aL24STGfxIvXRhNt3j34EUdyVUR5p2rYJWuE2H0/TSIGo4jg9z
6kC2lQzNBWibw649iCASWh+bL7i98s8rtyYdmTLujZS9/arquxvFkOFOkahoF9tWFdWnbpMys/Hw
9tCMrOZUFLFBXZxiJFh1VMjExVPUo/PBvZar8MMnu8W3S4z2NmegeF2X0DG6/b2u6uvokkf+zurK
B9Rgy6/tCELLAnTEBYqX11TioHPC/ZVoxhhDKXimpVqzmVaUyAss4FDzOpOH2uS+pjR0G8PmOnF5
L29d7vRWhNtwZCDwy296szsKxXL2QcU/yywHiLEG+GA0chK1HHwXSsi0RkgmJSDAOQ1GAHSPcqAL
oZHUPGokz7amoBUx7034QaelpZMiIuMo9KPzj+ps2AwST+S2YG2/N+/Mc+qq+xX+xBxIak74oF26
KoFcd333m+4FTTexIwds0ScaLoD/Df21Hza+NqhBevQe346HWsFOZvoS9ZUnExX2jTZkvi66jTVi
nehRQIlGgcWGzFUYcoU7l2FGvNlB/LDGwRTA0yBnRzdMSogV/L87TDo3Um2L7egc3iHK96Qr9RM7
qHHatJBzy2aczCdZ1Z8trLTz8sNXl3+xsg4y9zMKRUTrqpsZkDwBQWPWnHRarBmwHE4urtDdUbwn
3ZNuDeTYWEeXu9v9niMJpCGoEg9e+3sUa9/88VKeY9jhhn90d9c3blq/nhAmyXgz+WxjRm9/28Cf
FU7mwI4wMvbDJ4QZugWDxqSlcD1CfEEuxLO2mX62guBgZsLq2HAXoswbyhsFNGfuY/49rzoPpqOs
DJe+7DcR8iCjd4lxTmpFlZbvmeCwOB3wiOy7u98pVLnEofhzibjPF4UD+YPa6nNLKMyeTve2xMcz
pucSmzJEp8sTfcDetd5KA7nJq8ePnAez1BebP+87VNYujoxQEuK3DfWyypsFw+AdDDh8IBO6Qk2n
mQf7AJeJZVkFhMltrh+t6ZRu/0T0a0d/NVodk02Ze1+A5yLBR+ITrGdz1yhQUlP43kNEofVFNS1a
1lYARgYMNgEFB+nji+BwkKiQapRIUhQvHtDNpdjkldosOR+z/Wl/HaFhrKW3HlZTltNQP8oEG2sd
w9LK6RksHHzg6KGiY7HdvJjPsqPqbU+AxVFqwXwkuKNnOO0+4MpL7eRlcKlVZYdOjKFyUUX7Xmdy
O6xhiqEeZ0OBRt9cqqpWmv9tQR8Q9aZWasi93ZpF3JO9V1vMBinDFiBivkT96lB+zn0rBkSi90Fs
3AXjpxLHurDvP8Azr9bzJS9caeTEqfhaer4nYEKnufsmHjXLUuKlz1Hjfa0jOKJYLTEdPqd5TSrR
iMMutuQmJlBncj4g5FC7iJ8qFJX180tUtZMCJOKO6qXtb1rLJ3kCfM+yXk3Ws2kTfZOIrMy/ZBAd
MqQMjyvIAu0VrYGOxO68kqmIuJUr8r3BlZS1ghQysKfKGUQsh/L9neb2npp5A3GJqIKtczjyBGqq
3u5p5JLZxy96WXEIAFvopnnAPEP9R5udIe/JujJr6FYSsJgur/w6UD0FipSipUQ39WF8d2KswGvK
8lhQt/dIgZJ/UYqJo2xIkA6sjLAm9xTQ8QKhUNbMzXfCnewGe/FVqQo4ookHhELfd497qo3byI0A
7BI+2JQ9gQHkpyOQ+5I0hKbYk7buNMSlpnlXsOpyAFBlBEl0ojOvFxvRXVKVLBIZjfuwF9u3oL3m
cAwOZAQG6WEWOO4fdcG/8kgqA4J3chZoGsjTW47ekokR2Q0YhQCFrlWyqy33ooXxpxTOUAmxlvQJ
qbkAGadU23aadB4USs8mfyMsRvJ8LoLqTvZxVPXHXHHkp8ABe11u0jLABs+KKuDpsxRqDGWlkNvJ
ZReyvWvNi6AOCUKIaqTouRNV8gzqwamixa0e/P73w6EwdOtJYcun1fO0NgR3J9v1W+WaftdWuuOT
v8OBcDksm7p1mNNakEPUDP3opIzHXVTJ+G9cy0Ax0U4lmVQtIt5RrbUP+0xp6dD2a6TY6+BDO0c9
q83Gk7ckjqNSsBTBr9rNsdl/TYnFXxuOOvkH3AqzF8pOT4358+3lVndIzo3VyihiW2h1WRRiZjHN
Yf7asmz3hujPBNvD9HRNrXyfPPVZRXKzWM7JF26JA+jyY2FkzdSNKCi323SL2dKkQdb5QIJV5cC0
gnfl62sTIQf4m7LcVda/fjRTeE4PD2PCS8mkpwa997qSHZ9R6QvaWlj/vNKTwvvVPj3/Qz7+KmQ6
eFWM5Mc+X0e5RO0vzbvhJUBN0rokImF+ymcJk2MxRy7mhyIZoSwF8N4Ws6ieIqqSyWdmjKgAE/X9
IpVSHuQdpmI8UXAiokAz+zb49kOVNEMWcTaNMd0Bo+lJb2v6CJaLLWIanodYi4m3Ow5jJKfvPYyc
/IZCKUxcpJ+8idjDw9lpC388zzNq36jYCnX/ZGLvXqNJPLDR+ihLMDyK1ROW97iAZQpnWoCxbFUe
VXxLa0UWNHN3y1Mix9lZyuENUQw7b35nz01nPzcVCuRkj1XnPT9jOQKZNi4cyIcnCmbVRE6WfTQV
6WJ5Vimuj3AzLbBgDiRTkuE9hqSru/quPQvbJuKI18XGXcxkqdxBCDe/2oYhE+sR64bKZWG/AVPk
PuO7P3iMyMALnfnxt+SnXhrzHcQj1k7r6cI0xiKkAlW9t9X/+RpDsVePZo1mWyB0Xc3sSaVJPH8T
/wH1rwgnunx+GvZiZiICLTD7jQiVTdEdwWrvy5iWwRhvrv6kfv6TU8mfmKagrRox4hlqgtquO4nd
CKlLWvmfzqa66SnkDBwTko60u1eOQLGCu/xYl76WFaRw2nPXdoonQVBzxN86SDJyjyzlUMMl//Uk
RHcDF4o8ThFUUiEKfpyzKi5RaSDIoByES6BGy3JS7kIkw+TvM8ufNoPMnFSPS5QAcERtgJnc1h0s
Dt4bncsFpc/wnLpaID2jIO+iqnv7EeC/Xk6Iylj3D8SPF2R647zfKO2F2MwNUMiTLHZtSd2bE2GF
esNT1ZAPlM6IvGCX1MlfrQhOnF+J4VltA89jUd10SiWG+mQYrr6tUtRuZriCg3IbauEy30VXd9Oe
HhzWgBQZYoRKaiQL/00GD++auwtNYRiEniFjU7dlmRMzWRuf6DycrXBxvzkMbi97SNMqg6Jn71ER
2Wfly2cyJHX4yQwo+GmTmNojOuHjWhYMvvfnlWS3axhqwiRDdy5rc3ST692dPW9owGvPduIH2jn4
/ma2nWDy8DkBpZghHBTyBc98NeoWjLv/BfIA9iRrMNPLjioBvDn8MZA+X0fUVvKuVCvCPrzxaFlk
pR7CxYUcK7SF90OCsq7BAJHTZRN5m5ajpnXhogE0zF9pKsNYzxB64ywluW/DF68NItjRRjjtcgRl
KQpYITfaJMxO5/NUaievmEK+m5uO8suRpjWmtcH6Gg4XuEEJVbRltrZOMVl2gJiAsz3eWGmsDA7X
NvjlgpKc32gTGRx6G7HLp4ZJk/AHJAigZzY8C/+ay4aB8TvfP1Ima0DbaOmNI0rH8Ap/ZXkTSiBX
dMlihyG2NTCLiJps8EALlhVC5iE8LbcDDcV7WXT2GdHO9cOKXNAFamuWnIVaaHV8qD2BPESqRrZU
uQ7IgwR3Q1/tVN75E7wlW0FPc2Mnph6MNpePg2w4/oQR4KA9gCSrsG+EIiWVHg9IHJeldSR1zCLv
6NTAg6sWXt4O8VOfu4T27mcpGEFfi4JQ7JUhiQuSFqKll2S8AL124OV8nHqbGPg55xjvsn63ZoPs
0tLclVcP73LUVPQ7dS76kO9RDWhc0HQtDfb3mwB3YXqVUEkWY1yN0T5Z6+0dEDLqYl6VosoS3Ymr
XbmUuzil8+uMpt78Njm/AM3fQYXd0nqaGR/kCzrEljBSSXycl7Tfucz3s9s3hReRAxSsWf6ZLtve
TZokbmGRbzLlMRIBtt6Cz8WjbRk3bLyYsgtOAG0mUgYNOCr+fQWVHpvHmVleErWcJ5uOIRTE347/
yfkIn39PsH1ocSvh+AvrVbPkjeccgvT7yCUDB4eTohAJkkmGjGpjVO3iTKS9psD2iKlEAQKOjBU2
vbtSgiXJTO2IPIkHJFBUQzk3V9/pwP8Xg7jD+kzY3qFrHGtlix7ltI3jAxkJWFu3fextCJXoVBwV
ejxFTckG8HJBUKusYb3nBhJGmwbmiAKwFCJQIJB+LsYGmnFGY0zV4tXfbYKYxtcSBr0/RhHUSdMS
CPMIq6J3NBGbEDr5+wYImjEcX11Q4r8yvhk4oglpocK0+LmPZNQg4+jTUwKN8gZ06HsDTV6DRuI1
x1R55yK+sHRwNI/TWR0pEs7FcADk9hJ6I0sQGvosk5sBaN6BWkvroeA/JsYYZWcuB9pONnHTBoGs
dey7bMeCBtkq1S2YXT28omfLOekDibX/Lh4Fxl5re8ERnELMuOmJS19fM5rdp9zLw0AdEueAOkFL
auNmZNfjAC2VRlgZlVKXtDqn2pzHo5Nu7+IYlF7JbpYVOkf2NmrL3ZyCp+veqqFglyDGxSgnzByM
JgM8VG3PfQpv89pvwiRdke8V4opuW1UM4ftz6QjHlGy6dTXJKcnAA/5QbyrvMCT1NX1lANJrbyND
atBl/SrIHF59VTqvDzF3XaAk8cSE73NKa0xWnZlDqdPv1i79nFeAu/LfKd5mo4wSlebwcJKTkEAb
/wXJ6tYw/nMA9ZVPMMUPP8wts1VBGNHNVoWMFKscWln3wrDLH/hB+hztU8SQtNPvTqzbVBHdO2Rl
nc8b9LxId7MP3wxRtxVkx5LTGG0/T3yV8EISqb7nciJ5UVVsAWqKBazThTLiGE0tWrjCmT2ZSSoj
qREpUd1NhVTF7v+YB57RCO4ZGbyTaXNLAsmf/h4ZUWjXhoWcGVlG33XtP4Tu2uByKwt2tJCgL5dU
8j9qvJJxzV9Ku0eFRnRh8j1bSGvy5MLABvP0wnl1TQxkI7ARpH4/iIRsehj61HoDUQx/NGlzKxOe
JM9zCTRaN8G93N8JHJsySrWZxySgYyIcdUWOzdm/OpF6u8NZcD7zxJxyIEwyRH+RCPbPyR8bD6A4
yIKvKSDilz0ovKzrvFdepbT+jTZxpvUCIPtaqbfS3TyIcSlx+9QQW9qP1xc8LfWonUk0KJimOySH
6x60OBasuT4Sw3A5Ey49lku51BvFSMi6ntNVzuz+ORaH3GyWZt8ecPFsHUzJMZROzGPeolNWoovO
/EJed0AMikP5w5fuJOiJeat4S0zf66qXjMwA1aD7HQ2vnG9CrSCT6SYU8j60V9h+ICFvaQnwiT+p
M72dpD27LYQMhR9Sfkyc4jXv940A2q1YCzfOE1pLYd2f8OLPL5nL+Uf9WpYxXkDunlhd7w4nyBt3
bskgODB0OPBoG1VqpwZxMXVDx1ktUTkZ0gQtLQOKjocPHec0Yduu6gIUvIIfZybS5F5MK/RL9+0B
lYjAcsiYBHFt1ZLVumgJWaso5fhyuVpokrpoA/pU9t724Jg0N7dJETTVzAuXcb3UdXOvSTvewxj5
FA4n1+1cYZN9YWcYRq84c17FEAVrYm6z4inmZpYGZ2FJOUmpJQxsabhyn9PoLCT/Hdk2W/wiE6LJ
VSaneJvaZZkAQI3EI0oeCerkzFmcnj9Fych2vB7EJf2TbH3Ut0wpqa23yp2phnEVnQmUxfOzxZEL
TAxcwDvhBsAoDFWraoZ1pliWk6b0tPDeBPqVSb0RhlDu/DPgFj1W4RAR3vVXeRi4yyjYCER4XMUU
YmvTC6MmsqC1157uYfjQzdUf6jUJ1hZa2kbXX/CFb3LYyh7YZcOtpbwrsY+mhoer2kga5hDCSX90
+7d0gHDYx7ZaF9/Ke2MslrCiOg/jG14hwYatQ7G5ltO4+41LMfJyj+SNUeNi+ZEHdG9RjMoYX7Mj
tREFcFj3h11WNsaKlMEzRmY2yJS3WBByeTBWtqsACowNLuYc1l3doGHm0BKYmp7KoRg6iNMgv+5O
IcO6sUZodzJZg9ac2pUUWnwkdE8eaKyv+mwGXK+JczhaflFLeiUxjH4EZGmNhfRSh5dBRjBlpe2t
/gVmm5uyaEjCPcvFCdxhHra9SlmyvRb5hDQ/AqzC5MXC16AflcMAEIllRwD7ybtJg5G/pVpvZVU/
HbikFeueEdJVP/wI2J9FKC9QjX46Q/NTKtVlPaK2/ckxwL3wjeCZm5kcsZq2R82AzgiHCrJX+iYe
5rQ4/PKassQYksqNcjO6yqkdnA7dERZZKqnbmW0S0CN8KBtD1fY66Fw+ISTnOWesRgOFsOLzvZmo
uK0ZgpVwKQNS40laV5JQb73MoWuxvmZrcsLsLaaFBZNcSbthzhbfGhXAfflUzB6jbynR+gZI0baz
jhzaADjsGWgRA4HfNrzkNqNxAhzBB2wwWyou0xOQ0hJnW6nzVTsqb8rHOZZa8LNhzRqL8PCeKKKA
ogKCS6+ldEeLoUaaXf8qJBvvUqhnVQ5y2QfSwC6JCD9DILDv8lw+CwkMgyZgt5+pt1Bt6Rn+lc0W
Nn/K1IbS2Ml5u6PbdWzRXBMuD53rQZKzUJ89zcTygu3oaJCxoRsTPLXUbyRY9UkA7miMfxY1Kyjh
e9pExnVWw2u/443JZcGdBXkRxkTsLJxmFV6zTDir0thWmx4tMb13FONeWUjYq9gQshdEwpVVjBix
PDjoX55IhIpvWu/fp43QQ58/hwrSO9lCQ04Ob7mgGVzkwiON+whf5qW31xhtpd5CCQid+CH1IQOa
g0DLj2Osju9pR2SHQ50YR4EI2xX2G9kgkyXl3n2oZ/QhhZrns1lXPD6BaPayXrkn6QbwUt6nkKcE
ujtSmJ3jX3gJga+F0XMdqUUiUH+kY/U73m3c7PTiiGgUq3jJkVo4N6w6sVJyt8iyNXdqJkjEMbjZ
ydiyg1JFoEAinge60ttNtZ0IsBbKg7RjRuM8IP0l5h40MYEhCH1Bu6BG94uo+5FTaOjx9es20NgA
V1z9EXkgyV0VKE1ZK2v3eZ+Z+UXbIbSA13vNq9kiTBu6+2QiIIvmbMo1zAfqYx/IsKe8T56TfjOQ
woorktbMhzDe9FeK9CAVWjTxSo7ddcnjiNcP731BTv9k74tsYEjM0v1EobHnLKs71+kpZhDutCtF
CI/c1ORle+cS2ZarD972ktkbXyo1ZwjIqoauIgJy2FSMMr5fOi4CroZ4rC+iCCzexB2l9oxZKQfr
/OAGNs/SP1Dn0YuP3mhtHV8b1bDd23qDvw1SYj/tBUollkuzUp4+a59Yi4t35Wz7Y4BC29Z9vbhx
dZ3WUbSnse3aaf2mRmELmWEPa+nBIxasRm1EtlT1+3a5nH5kZQD6juHbIU+R/mfndYswHNr98w5p
JTo3BovdxO/2GR87A/ZVdIurRA2qm4rCIrzh2gpk/WvQzXEmDE3/CPOzYg94idyXG1Ow3ybkcBM4
U1mexVJUNpQc3mS6uZ5nJCtV9REo71izxSkGmFW+puGBQ11x5LiqqIwAIlvjKasJtH8NnptM/VEt
oMe6ngfKE44+e5aT6VP7fn4ObBTS0UNg+PIFbCMvVu2RALrKDwyLPlLL4TrzwBtDxSgZmEJmxWGq
TwC5xkYAh62hHrwWQ3c3pVa9mAHLuc/dC40argFit30yodQ5xBUSostnmH8KIVDgwXARL8dmljH5
WJX5NQGjl8uM18B7JaZUn9ExtUQ6sk5t+10FPZH4yfa5Q3Oduwzk2NoeIqGlX7ROovang/5EJNUr
jSZ92wyxjdzwHID4vUrjUdfj/vBL3DBJ5BER43SJ8N99ePzEdS3LTByT+N/ntLsGKNtvZyNBfRLJ
dtR3Nxj2xnc3dbsSLh+QTDYaKgPCIsx7fDAspaMWVM7y2saPGdgRs47gq7MPTR20zXTE1bBLXOwU
i0MwA0yOL8BT/PAN5JPHq7etgtjUmykx3/lwvLdLVpIh+Uy+dpuNJ2poyz1deBrYLtV9fVUQoGr0
dFQFs9q6WKOmQ8DIwDZX17XPSAzTgBfxe/qK7hWT53t28b7Ajo4UruQesiThPvSnhmgWBcNOzfQf
YNTTJaKAE+Q+XtbK5t3XcgCTUptPPt2tfFQpx22V5p3gzdaGoADDUbWMbqPKmXvDFDLZj1G6S3ZZ
LwH2paOysTPipuJeU32fMmc7Ifs309y+81fRlUrMt7EPPG0FtMrIoYL0n1mqfvKIfO8qgCVoHo8O
KOWFPrzsy6qSHCetRlXAvqAH1sR46QKxq3peLkiDk6DvxbMdToNPKkRyOdZJrL8eKsXxckxI+8Wl
HBwhrqSqcRNDEM2ZLqeqmko/stVz1ysUklboYpUsjVEVHwLJUXH/1SBEQ517HFqXOXLg+QiP/40l
DE6i6CcUp9Dwg+3zciCOLhU7TLANtyJ7hr/vJW+o+sXvXw5PG8vQUq476WcERWFAZr23KbACQcuD
L78ZBENBiLm6stdmutiKvdwMsccQuYwjZ3WmTZafT6tZAhjnG9h83H/PyioorKoJu/PK3IVBgh7o
wDoD9G44aCnFm5PGF0CdNr+re8z0wYETK/n23i1GZs+zzqJ2896TEqzKH777ttJ/D/vrYkxtbbUE
il0VJaS078+G9IoZWS5Xwv1qtdDFUhUHNaMnbIBf4Wxr/wLyi7qqIdNSMEVidMev1RIUENSbYih1
8pRThcVRCjXRudLCsk8r1Lzag3PvMFwNDe15pNr+i9HxMg9wsX+ksae7alR/RiEvvgEsUrCWmrUx
h8FeZ9dE1Opzy+Kd7GrThJwnfZ1LLYR4htjrebGmAnt5FtHqHbqRhVo2vQgn+gRjYJQZrv2mYA2V
Pt2cpJBJRzzDMGc+zmMTs3Nfr53O7gm3pygNKfpJWNxn68rFcPhScoiie3kNwS04V4BN9izuP5Wd
OWWqwps8oIqaR/K/FTNA+FeFvBIMCcxboS8I9cHHgGmMfc0Jg160pfIFeVE74LC02yDGENi458td
gSdLM1gFqK6tP/dsJRqgU27syumw94gDudnKT9n/KTcR9AFyOSr2Nq//g7ehe/u7zgBWtMCQPyJp
yvaofYAZw7b4/LmIIGVGjvJHM2wJj/ACpSdrpHb0f04wz5010DoJbfbbdv7k75yLaBuOcCNsYLqB
rO5cx4s8rZMC10SdZWc3ejCt4EsKDd++TRmu3H44HP1HAgyBeAtVMWUOKAippwS8GjMRYwES4YJu
daoqKaLGWOCpIciB0ObcwEyiXfm/PPV3ikkxIg6RbCA8himFSRA3D36Wy4nSjG/BiXSLREZO8CEs
jcjAgt5LIsRW7EI2TwtlaNK5XA1jVo3toJlvg47BcA0Tm2jUbyVMNYyQVlnV9qCZX3gECKey6/rN
9agm5kbbPLNt3lHBUeRz58V9kg1+pFCfmjI8qMv74ZrZVy3bpkroo/1aTcOzqLYkRXB2CAObrm/c
GGMjLhcD2nV0N5BKt301gSh+g3Y97CVOO1UOVykuIxbUyRbfsXOBTuT8dSeF8rcYraxx3ZFGVw9m
dxzRNxRyDIt5KFfzZ4fIavlt7mPjau1YbgZCvKLFahJFixpNnDAzo2wzbLwE/YxUPLl7PSQCKgSt
t1Oue5ihmx8JMVyNQdKojTa/dLfM5jKQxCOhrY8gu4of8GjND8OOeGcC6cMXSFZs+pYEjq91kOP4
En9sisEitjh8Fuco4oZ7qjLN258YWeBDJTewqp1q5AGbYvlmxsQM3p95A07Hv72eEx3/fARdN+yD
WOIc3U6XG5VbyzRBEDeQYXQQE318B7Xd+2r+Z3Xg1Ns9U3cv/y/hS+LmvqzwanjP9wNfK8tHbQ3r
HAxMTEkpy5O+8ZGnssiLFdsZSjmcM/5v2LkYsX2xYYO2IjYpU8Y0Uds+MCjLimaBydGZ2KljVtVS
yzT083pmefNtBEx1J8m7QKGLlQHlB143pF9mkZ8g//EkbT/L94yI5/+ov+k19/jPmGDHf3fWOHHO
J8tPh+lD4TqR4BBb8+QxoV0MjGZSQ6pXwGLs9YQwwetw61lWnYAqLwUUzE7L3brbaE/FvJgKyiUJ
pwKf+ndU4kdei/ZcwZtVmmK7xYR4EGMLGr7lg2XLfqTTqSEjSgNlbdSkHKFvhxRCbaZURSXkY7XP
9HLa4kC8Riv0aD0QmBGP3xlS4mePSJ+62ivf5QpoV34iyoLy+3AXBGHHH8txNsDuJY52Nc/i8rf6
NSoNCGXyu+XcJpgULJyhzpB864joKp4vPbUOqXWMLHK3C1xi36ciAoqOJzVMom1X2lff335zanT3
oC2Fs7eb3wHMoEt2386Ba58J1RkEk6FuC+eS93rMpeO7eHFLX2huiblE51ld1oHw67iAvRyp+1BQ
ZroirSE/vbjECUonAyhwPc0fdZnc2VVy2MNbUh80qLa+FH/MNl793g37RSEd9ujU1lwFDPF9UH8q
QpQNzUz2KxtisHIGPGMRGafmS5MLnZQtzgzOEbqCtwrlIkU0kCWZf6O+PF9gJpkPiM7Jvri+/Awy
Wht1wVR4+dg9WeZ/yAGQb1cgvAHqvcHMh8QXL9MVhARiZhwJq3sRKYA5hremN9Dg3BofPAMuPr5w
wyyoMlEBRJm1hCSe6PmvJ1F9YKHtQL5AfpBWDJjd6RNVqKzfIar90qUJRpufYeEITcxePopGE4ty
khVyUXnz/xUIjjMfqFfUlzbALwf4pFtLTlj7vSEhx8BStPzUgrvzDuGUTXnLpLwmaVyxc/K0ZoDj
3JWy0rRdbnogyDgtan029tHImDRhWFvd2GO2Ij1IkiaUIxG3OFuGIfIGppsA+OZymUpNXgLPJH+X
IwuP2/d8GTFNgDqmRJfHJxubE1tSm49qebFsTKMZNRJcCAVsrHIe2pTE69vT+qZP21ZWMKdA5vHf
6oxfrbcC6LU3k3Hk9MwnVhZ+oTGFcyojwYa21Eo+GaiuFmwAnRKNJFoUdG8lHuxBUsCS1RJHmucb
cn/8m9CVMHJikK0SSL4zV8UwISBx2NOZhhMlq8ROipbgXhA1vfTOCaHmT/QAQRyps9tNtVYilAUV
yjuUiAEhEGWNUAy3Eo5kwH3sLd2Z6F9AKS2mDlJcz/fIcVec7DuTNWgQ6in7ILJaEIxOFtwGAbBh
pxdGAiorAFZJKmq2uItXRix3ZxK9yeuVxqaeQUJ1IdGcRaVkfH8lUHJVQ7c8QfQpLuOv4uJouy8V
X6aj10t2yijiAKfdeIZBF9BR5K1jNyaiXH5OcSSvo8xmZOvQassjvE/K5gZVPE/K+1o74SFmgVAX
p4tU5HjAfu5OQHTBvV3ryum7L5iED9oYn+BPpgBNORS2yFvSfFzae8EI5CEn/mU6cfnQlpVmsw3A
QHimoByRvNEpl4YNUH689Cn50h75IHLRolwDyqTpdLCM1vt+8mktRn3xXNJQ3jcICsdpU9FW4DKu
RuE68jhVOfz7u44HY+xIiA1EOIbuqjkEGQoup8JfMEEpDthZk3enZTuc3O3qUKyAeFZ94fSUwKJQ
atQLTspnQTj0FYB9FlIhbZS0neFiiGCrTdErWqoQQfvwPDyN8RrfHOkHu6NrK+8+sO0Ozy07zBrG
d7FA7IMxGxshbnmq4GXiJEROd1W+8E6xq8pjXIe3Si74UzzEloy66tSnu5NkI6bcIbKokSEv8sj2
WeUUyZEIGICeTDS0+E5oe2npokfIzcA4CdZ/rV1dTG3G912D/PEH7Iab9KJO10l/h1pVYKdcB8R5
T7YFrsZ7fyUIcGzI4+iaqSBzJ0JguNOhIyq+b9Zv41YxCbnuUN2eolwbnUpYk4urOEEnI1xHJx87
a7QzVUxTOPjhGXuxMItbgswXSnHstoHLiJJbj7/guiUtOWdZPMEmEGsReL0JD9WzSzAjH7YgiBUc
ml2bpqPc5tqhxxyGQq0OFbK3M74yKmSFEWZO8mZX5R4J8yg6puw+atptGI2w0qumKn2Is+QdOU2p
qPaZqWCOx/xu6ki6BsN1RUryWQtm6aKd2Y3Ir+G+4w/+mjiqzXzgRs/RfU6ZgiAsfhdJUoNdlRhG
z+EHA20jc/tFhkzKruyj1ryEFP15+96p4GntLXv5yFSJ68lSGYZGGqdBkyhDnldVPZUMRzWHW0eD
oYWYMbxBCsGN4s8i3thktfa/bxXCxkchcT9O7xT7AP2CB3ExvPfEK8JBzEaIE7TZEulBPaNvKqyR
AQcLd6lKVIeYt1XZcC6sOe5kEmaBaIyXZHswmvLzyVq+1ljXF0+gMgHGE5gM7oee8eXFgG0CevSx
MC449DCXgVKe8YjT5YJ8gz5LA21s88EKs1M7b9Dym4Qm6CHwgLSIZSZ3h8tzhSfn6Bx483yjXJTj
wRPPC4lNfTHkDZFB6bWOjHjW1hWD2sfNZy4k/HJKKW274K63X+xkWdw2xzstNe33xiEjoRoA9PEk
9v6d5W53jjLMESOqkjAnxWcgP3RUwFQeL34wWLFXN4CkHgHUL/sk7mKDVB/1+NMEi57eK2z1Ltjt
ytWPU7jULbGttYciw7lnCQ6BFDKoil7Or2ZI+NpAnpKR4VWjNmMvh+dSpPRtKWx0SIHY5sv0y+lT
jhaU2cI7f5lJM5v9SY5c1r4npgGTz0NdhmrABZWrQMwri6Z6vJNHExgpv7h1GwOLuHzko/V8TIeE
FdCLsAJtkfAMq4cQ2OIaCz5T3TmnST6c6ttkzCrizcriNCuil0H/W0AacRCEQGqXZVTsPPi0RWGU
vp3HeZRuzXEhIty43yNoX0m/UK52HT0ooDw7DOMDNrZI4F+kDg57M2i8QQqxz6xWZDFhnIQ2xsT5
ee6x9oSAuedpZhc4EgLNqpR7IOkrfv8maumxaRe+mpMCoXHuG/WV700eRyRitahkuUu5EDBZwt5F
WGK8WTPcJI81WBI0V9EVfZWI4eLw24u0LAJhMWKIU6/hZZjOlcakgjW6KpJMJbfWMT2Gh5sfMWno
/IicUoEpLZTtE5lJLVckflSywQLWSgXwwoJgtq62iosh4pWeDO+QVFPQ5jYIQcHt3T5E9h21eRjU
NWzEnQPKcyn/FVY2Qvu0EfEn9dV+5AVb8GjnTRqsxfpeuDlnBHvnBVJSZ4jmyw9vbqe8bC5bGt7k
SGOFvoT/VWzfCEl5X1JZD6i9ktcde8qwnwwqpEnDX7hra+g6TbYEMomov6LBOLn/OKaQi/hLUsBh
RdladXMuv7Ts2itLctkZ+mCRi4F3fj+zHG5gvRseAgKg7HBbk1bVNUC4uKMewt2/Y1Dp4MZPUL5W
7qkx/9IUjsB3f4l450G2p7edRd2TzueTR9Uc1ug5QnTi3zfZu2DaS9UOigDcSB9GpFnyaUKhRsRd
OPcea5OfqcXMmAuitDYfNyiJGPfw2p4LDSosUj4T5XnO6yGYIkN1A9W8N1Wrx7qZhrjirCiOjtbA
NTgUXtM/kmiID3U+ZjkZBnS7fhPB2aGJAfOXzEvjcVajbc4mBsag3wLcUbukEkzei+FPVuJ3J3vS
iD+RUC4Go129PmWAONkdl7XJU8wZMrErIaiiNEj4egU+mPqzUrHJbe3dASQOz1oqVc57qydtDokc
Ws5CZs249BczRSKZAjFmIHJa3suncU81luluYtUq5fgi6kLfHwemk0j0F7eV5p8HFKUr+/Ah5P4m
o9bejVxZSPsazfngcuz6XjmdSE9UENMr3PFOw9XkxcO3U2GnozbAbTrE++4sdcNtqLBLuzOWZtzy
neWzfWThvznS54xjOQ3ZkJmHZP9MCL/pSCn2/avmLQ8O18n5hqB5DBLL72TpWl1E/bzyRXC2tguV
Je8IwJ0ePRNplvB7AUUmNnAgGQqwVCBuAZyiliEo1/rOes7uMCw/kYvApKIO9SkDi6um9zPMQZOT
snN87CV7r8RuwkIFYM+xg3yXKucCNCU7jajNsJ4wLMobWV+IdpZ7ze6D1Dph5taGEr2ZZ50Ov2ux
oQF36GdPh/u/TY3hihPSOlm47ujx3rU5Da9I9gK/WvWCUIMA/Yw5NoBZjLQnwc1dnt8W0HtBGxVl
msepL21CFanh28HYfwRDlOmVknUmixzpNJ7I4PVF/0aotzgyO5g3cPj8xDnF4x6s+w6TU1O93eAI
7ixv9+g/4MO2DRycScLPQ1ZsDa2gZ/SEthgX+YbAAJUdNUsZkBxPLJRQvsicCHTSfC5q7UYcFYn3
23+KFUqT1+kGw9Y/EvqrUf5DfD56FWPLxJ//o6kgWXCeRkyXqgDsbCMZ2oIYFSXpYeLoZrOjBQ62
c1U5DRk0G6hLuSdr3CnCFaxvbzGJPokxl/xd+4zGAA3BuQj5NQxsc0Rtn0jnCBaNAtUwXDnOJx8/
Kr+1I3W2TvU9AkQMuoSxl9Ctm21WZmlKe0wlrCrZ7e6rIUIeEN+6qDJIL2E2DXz62OP8eyw9wfgx
YU98TJZfcFnl+gPs6T+sV148RPA9Hx/+hjl5CYQxfu37COUjn4t604f82+0A/8qTQXgEShiMqWzp
5JZMjsyQHuA3WcX83QgM2po6YE9pqrQezwiqYnNLEpYHugbUGoEkTduT17nexFhxcGXjp2Y4ZYUM
Z9FjM5FahDdw1VYx3zHp4wZ7FSh29sXAZ5KE92BhAoH2tRuRcv7fRTDwYUim7x2i41nTcydSrqxb
ThjCFyWasWaMw9n9xLHotsmDk2b0IXLNe/1g8SRATFo6OSEF2NawGKfqBv6OdsH/ErQRnXKoaVy/
omhJJ2Kv68Skjq/vpLlMR1/OitC2d0JKI8C1z5WeCCNfQx1uVMu7vRaZoFfmffL/f/9eI+9hrgQL
uGEPTvBequo6Ruy93K0k8y/KSh6bfKR/2sRlOyTxEh7qb/wMLbA/fKyi6KuZqiHH8akpkv/aqsM+
GZnI9iYosOUG85IqU04r/71WpVf45dYY8Ey5H7GSKtainYYNBxFASoVT/v2oY4nncsIv7aPNgCKj
2xFluQhgylEmpYLJhKLXRvtgrVJDIPS6zqXwHjCoD6olWkpnJmAxKdzJcl/hoA8JZvdnu7tl72Zy
6TfVc0ebnN/MGRpAwdQ8sqCeVmzv1vrBvNbIObbGYzqOSNSEruzACB5B9RIBB5x7gy+PWw+0gT8/
9zMOS7cwyubHNrytQ9mCvTg8PYW4l9O0b2Anm6dYfMoNnapNyOlH+6H5PHDdf0/MeV7Mim9v1hV7
71d1ZlhMMwzFoXVVzSRuYo4TCMhwAQQWhvCmyQi2ISkyknLDrSy7hf++DU+ChTczq9kYGG5qSYHM
Ofcr//sy/mT3LA7vrl/gBM/SGKN+8eOVPgGVonusAodSqbp06hduOpduOjMeUW92BWgyYPV8CGV0
vjtA5cyUhU55dzxQ6mJnjJ8m0ETbB4biOM0f1CW7yuDA6w7eyScTPW+N0We3R6J4Wc8xCRP/HWCu
7r17xMlO9EQBzNub/4TT4+kPyMBn8EeD+H7j77GfZKYXKCG9OEKQighxrsl4rb4z3DSqnC22AE+L
4Bg5UtHBtMjF9r6qvUVaOypYrQRgKJZUDGIhvkaZVth5Chajm+H3MNzI8emDdQoIF9tvrHBjMlh/
+z5arANl8NXb3xHt/NquV+4HtA21HSBzLW6qjmKlH18rdKxC604CzdJvrJo7YlsZDFIkzl91nBkx
XzqcY4+m6i5aj5fwkduNH6YViSIDp0bAxEAPb7L6NSWfQOWLbMxVhEVQLaxi6wJZuxVvxHKHb+Dn
FJe2iunR8qQowxBWCniUftoBbm1ntzET6adrt95NBPdTISBGHBRCqywAOj3D2rKqY/beoCDE4b7i
9PbEK1Z6QEReQzm41i1KL16CINMIBpRyCPbwZiObPzIrPp0xJC+1CFDwgxzNLWkLCixxLz85dPsa
r9X8gN9Vk2oJ5q3L7YPGgZLPe4B+2CGpNes6cNueaK5JxEeyqnpPooyDp1LQ575isb5WL6XPyxAd
D/M/hhRM96F4HRlRleyDzij6gVvyeNwdrOp9Upz2qLECXxk0ILstTmQ8pPVtyhO7UFcHV59WDiDU
fn/zOPcLQO4WWMVYm2HFC85Y+hwAhYjRNLX1r6J7QaRPUv07r0K6ct/TcMlxUBAtexA8ouo0VrrS
261XdVEaM07WktpU5AuJdwUN9QV6ooEWmVF7xPWH3BmadRsMrDRt6FyXAKuE4Tyee976Rlr8wuXc
cPeA5SfFUCXChOzSljNKBHcDt3ikMhjZwy2lBzYh22VKCmBy6kXBRvCOh28g6T7fCLpDmzYcl72p
vytMjqW7oxxENwlwerQ3Lb2JSCN7ufkDPlh2l/rWqNMM3Byv5JYOfEfSNGv9hroIpqsD7iX5hV8e
3ui0h3i17lgh8J3NhRVQpuGThXvvmu5TMnoe+I6nxGoz0tzfdBYLp6pHXOirqCFzJxKM4AJuzAEa
2fgVZNUdWhlRxf9SoUYcv8QoC1OM1vKz1EsUprwCZlKJV1ihD4AsgggN2p/L7R5FWgUe4vf5a1qN
JvcVupSHVuOC3ibVYc3Id74qNXwqsPB22xrIZySka8USsuMGnaYpU3UnOiW/xHLvtj4ZvecFsIYw
wBsQLilAWMP8QbWFt/9TskA4P9SN+ztztlVzj/tChoxZ3tKhYrgNN2y3P/rX7ZaWF42V5/VhCZ/y
ad2vxRoCwx5f7HeW0Qu8VknC1rWGEEH0rV/sh64OA/TKlxc1mwOU9GCDNuXIlMCIRNi13Qs8bSD/
m56y6pSa2s/EomwwD9pa2BhOx6vRj9RWdOTCG8Ea0xUUOfofAF41Nzp8xlhDf6Fr6p5DJliEDyA1
5A8X5WeTmT0ARIZoChGtyBpR0KlJ04fGY3CSqZ3qeEy6/uELxIhTaAnuTRafZFg5y+OJhTPLoCDk
HblJR9OA6CCbr0DbgvOuvLpbODwpXeS97jBnHkaToBoLPmUKzD86R/zFLIHWeSzuLYNYczCh4Hvi
MB/Jr4cOz6WUEGXzkO+Iui+v4FZzVYfOrbE94s+Tu7Nn4WB9bUZ6CSzCu0pzXaIx25qckZE/p/mA
+5/QOwg9ioweRGzml+p4VKzC1Nq51MKVjJ+AOk8QWCXUQZzTCXjxlR4YqYDxW4XNqTMhf14fKKLr
3CBXPMj7qZPqr84cAGIdisc2lPeUoJayW/6rzcNbO7rQ09dDOH7SHRRxfzJ0uCmv3fCkxIaigWLz
W1ONXZqJeDk1gaAbkDNfeRZRs6fpOBg9czPp1ICerh1tIUcoAuakVsXofURiu5JP9JIKHPDpjoYZ
HhtZOnOVSb88fFN+1QTtqfszeaECo/2xG12fyEg7nh+lI6mSivQ/glCo6+zBOi3O0aRlIzeorJlK
aofpFjSbYzbGOc79zSD+iCZwfp5BYPd9el+4v7FFCZSpm6iWcXTZxWArtaDXnYFN2BW2WW628CAk
hUB8awKtZq8e/fZb4C39A+jZ0LDs6uR/AC6lKzwA0G0nKrkyrn+Qa+khj7RiQmnDVquxv2u9ekqH
/PsPwS4ve+OpqoKY69RyzlKP/pU8w00CUuQV9Gol9SD7TySVreeLHkZFnsiNBsVbZgfNLkmTp2ly
mKewqp798crKFcEs19dTodqBaFExEf0kGbh68rDZHiQRa6RVjuoKHuZab8SIiuX8k+hJSdeCVD4E
zW+pYmNqeRMM5ZJhXGKSXAVzAndo8l7bAGwsrk1HC4Od+gOMeQeHVZKIveX3X1jPjW/j2JrnlGeS
BacK4YgMDPwr28Br9hKaDLLo+YFaz4z22KMGTM+ea7poVIpCc8TouomZ+PSySKYWiQmVZODWlR2v
mquWgmhsFxXPUMaMqkvIqxA195X4e5ZYh4Vhk07cpd4M1Fs/mFSmQqXpqGfuhr4awdTHBK6wB/in
fST0iMRah9wTUslt8q/DgusZuBT3TPfTFDxsv7uxZTrU4my/jk/60goePT9sFZV6cQt8NDd9MH/Q
z4wOYj+HHI4VOyt75xWBDZEA0vGZgvQCvMQX5Pq53OQDYkh6Uq/gbqGLwUXfNZuu5tf4yJvGQWQE
wNvAGBzvwD9mjyjHpAE8ASOXN7on58ARQI2ly505rqUdRqnnoBcgtSAESIuzrizLFlnG1bEvWIJr
0OqBv5ugrt1IzQ5JiPFPgC65raORP0xCNrXOXiDQj+gAWTfXduLT/Hmvr+YmNiz7P+i30AtRL82N
XHco6DpaW6cfxNGAw8uoq8lj6Id1x7Ikc2y1ub/dZT10J7mQt88gZek3KRtX7BtfShSYlBgerLHw
5it1AMnevI3/qHecA1XaZksTPn3BqL5MR63F2kOHx7EpZe8jKe19klNKMIjbwruDyb6rtnYWtLeI
XKdEq2VSe3nBHyMustiLJhR/w/EkWhfcOIfAOLBLmo+vfPVoxcRoT6WU8n6KwRdlKr60chrJco5x
de4Zxh2FjRp6X+Flb9+NN3AcK0PPQTwHLQP8DjtOz8yUoecQz9EIkJ5CexsTLGTK90glH3+8GpYK
nrdYJXrkGqlEKQsI7IbhN8tSZdXL34ekwz9IrO5aqETF4SGQQv2Xs4J1XKTnL3PkMwf//qCCbYAi
TAU0BtcVzA6lDdwkV1oVBqr4wNSjgooKhm2wsYFXMgBR/ZMeJmsiipRTUluxOlkib6JXCzZS7A8s
FZKrIoaoCiUvK6kJLUjO/hKGaca6oiGlehNtUsvKfRKlYTv/2hAvXiCrs0XXFKOnhKkMIMSuPX/o
PlABL0HCnCJYFhs325+d5SuPhiFQ/9jub2TMqfkGfK9FZQEgIfTZ2IIB4z6upcwrAs1i0H0hplsA
SGbxvtGklMyIKen2eUf6uRTwM5TxbEG9sXs7ZPGiP+Y1ZUWGpR3LieLgx1MH6vO4Kapgm0w/J7O3
6f5M3BF3mzbq3IV4lJWcGKMIZ4nvgtfoEvzd8nmUPPy58H7W38htS1/tOXvFkiK5/NcuZsj2AdRC
NchKZdKkRVfMpJ14286ynRuqg5vfdn5C9jlIXhe4OaMNW4EXJDlWeDcgPsb5rI0fu0tbMNDLrc1o
aIMNAfO6GMM8Oi7AibgiCcSNaENltKqNMpr9BmoE7PJQYar/gkz+pI1BMCneZXaoVqayXjuhKxzX
Fm4g5515qSv1zYF2CHItMpnzhCtZkdHIZpUy/O0FV9iOz6dumV7Jrt0JbccB40vfWl3clCttf6Is
usNmZSODQfTOiK6av0w89gPYeIUYgbWInArr5sV2EGbzxFNznvg/7F8MKMJGTkMkDCoAxLHBA2/j
yc7fH7E2FEV5d4JlAfokV2fXZ2D2Jb/iVrjyI0yfpYACmzv6YfB88ouCNY+adP9iws4fFJFTZ8D/
EjFE8vsMcKzwrW4M/m+wXzOIWUAE+YrAUVQUJYEawoCLTeilDDHg9J0klDFxIruLD64s7eGa7P1H
kuDGA91TDR9UBaNV7tsuXpuFCch8Ou2OS5vmdzHq9gLLe5G7ExzYIWxoSn9imxxxarH8FXCYm+ps
ROP7NZ7IDhEJM/IEI56v8R9tr4ycKoiVTKNwTphcDpaHk4hu5+ZUDgonnmqp51IzPMcbgAAJE3mb
Fe6JFL/K8XLej1UO6qlUAVmLwxiyZ2XZ8PcdlEwCxnk6T/aG+1N73uWy4PV2JRSawqXk/RpyGog/
eIURuYaEEI4v0CcDtgIqfhLhI1ultq2fyy6Ks0rCbpWbz1YkLdw0mCmXvKOIE/cJSk5UgKqcV2Cy
DZJH9AACB/FRnD+vJnXr71+8/XWuZLzR00KnasXgxa+WZQ6zS6TNuk7OZ62z2Pr2/VEqZBvJ6gQM
Kx4hFzKCfDOpP3DfhNIOZsycnRoNoKJcGCpy+n+fqP9ag5BI8A6k1K+7Eu+PMJvfHBHIJ6o7MPsi
2DW688Db9srPRnk2HazwlTo9dWTc7Gdeqk3dW70abu3Vf5jH6TQzPm8n0uGHqow66EIKuiXDkJuh
MJS075LWlpBscYn8OKhx92BzN3Pu3qYHZF4nRwm60ZQ0pZYi0ruZmZi/BLaTuU7FM8CwD+d1MNaQ
b6+YGs84JwBqKqx+ui/LHbfIqGUofFK6zUBjNHAIfknxkyJ2P20tWVafnDITMbi+4g+o5g38ndir
1COnUO4EKmy3zigJlSlF5Cua4O8ec/OBemL5pjpReYEw/ARNC9PxHQeEPKj+yPPzS4WVu1s94MDB
AWS6BSoaTjvc/u0tUXg/jPBgXxXISsZtuQ7ZO3LwwEBSpEuqZJzD96duT3M0sOC3TAWyWp3JEDEr
ua18VVMdVA/1tJFVV0IIuE5J9v5rzf6tvuuZ8eGp0vYxbHtrZJf8Y8YvXNM0qLp1vSlxu5mI180W
BNXQi+icFzNce/Fu4XcfpGT8W7QSM66AWBCNIBDobojfsupEzn6d+NSJkVsHWKPiQ4t5XeQ9lbmH
ImrFCugGEUEpcss7UcXK/xEpShJAO/Gd0eBzsaCr+yeFgov5jq3/JQLXZ7jH6Nio6TNKbRaMvk26
xf7QIh88s5Hg9qNQdLBiQVB3w6QLRln75VS4gwb+Tt2Mg/LRC6Pa+D3FAtLilo99JmeiBGLRZXqF
5fD5pfbbqlSTcqoWlJR19jIoqh9VH06ec37T5VZ586ePRLf6mHtVy6zH/v4TDrkmNRO4xn8dUNo9
Ed0a9/kdurcJV1bZ1Z7OT2Y5MrdZXG+PuWHzdq9QXAP6NKYwH8ktJd3ZDexB/zeou/GkJmUMT5tx
v2JHg0yKuT0N0KOFD0l82Urv+9L82XrFtawW48bhLilGi6J47v+Cw0nuFsBRDnsk7XBo4h+2UiZX
Pz2nbIApU+mXqL0Ta8KJk9EQlLhTP9CK213S6qKxQzJVxWaYaITX/jREeoLok12EVizzhZaP/w0i
cMjIpuJAiowt5xcuH9buh6eaaZDEkCSlRd7vZ572jEI3iDrjSlfXTFtZzWOZKiOJBAQ3PvJWYcc+
9RN8UYFkIqmWdBGcLQM026+L5hkE++rOkTgrwW1+jn57Hs2NsS9iFaPjXBX75aj4zHR6+4ZbLyJC
LjfZy448R/zAPOoqBRPBSKxv+rM5CaMESdOYH2kbBgbMbuzICLswB4EHA7M6QpjXkjUF+iof/dKQ
0awaZnOmWhntAx3PrBAPiCgclobefgA+ZDDNniAwrJmXxvP40OKq7Ec+xF6xdUpV9G088jV+v5Xu
9Q49t/XVI9Yc00Ni8/hNCxVDTFErIrvvz3QnXgwbFHPpZFIo1jh2jXLM3f4+knFjDqpJUdC/UNdt
H7P4WN92O7Qmqwhlw1WZNRh2XZYaSiERDO1q5FTTJG9vtutxcjHb4fHGXcbS0QYbQmgmq0fTfhiQ
xhmdqv5wKqx0v6lWt4iMnPJv4L+2Hio5SckKJyjrglnveVati5oLa37ylputsufzPJOZNBAPcNfF
O1annawKVbpprP/y1j8SZQGiMG9+WxFUdefk2JOQPMz9WEXR52GLSlgHh2Os/83SrYAv+/cq1KnI
WbPflulPWNKbDMAslXIIryFI48GYHE6jFkcn+E2iHAMMuD/Vr+03by+y/QfhMKDp+GC28T2ZIPuF
LwMDlID6iNfa5ohJHaUeqlO/+djUxGU+rP3O9gp9wAybwK5O12mgwLeojSSKHKLDytxdlvRIs25h
iHLVrAiAVVBl/15KBxvfXmkQvmXP1nVOwwJ9H/cOEehI99FOtpQsbc8XpbjeopSxnlak1PEC5SA7
C5ugHhYthS9kZns6C0hOQ3r6Q9pgN4NR5fKpqGyhBS+r3Dkq58P2P/XVz6aGHAmnNrFcRJo4FGIH
Me4N+cbqbSLP3Dj7jWVpRazsWUBmVivgLDaPHA9XAKMoWumumB9PbCM2m43WWZT0i/qdCnhSAtt8
+qPBXBIP/ZB+9v6dCkccPyAwVoNAaQcccQnBC+0DWHcsBLORPGrUOfX0vVV1rfQNCgRT8SIWyqPW
4WPyf2Wq8U8Y8Pz68xFtll7wK2YJO3q8TIk2de0KgyjxBBRpNarDla2L0HhNGhDTSapvb0r5MgTE
FDZ8zmwHZ8+P6Kt/5PNmkNVDq9W4kU7jira5eAXAMVR+4WIDLMhbBGWV4JU1g1q/3v6BYEL+9Ur9
yP9psD6VdIS0eSWjEn+3At6YAXVjry18KcC44mRLMxE/tODqxVe6gAm2bxAEb5v2Xbv1jWP2Bf3Z
oTQIehF/VvtyHOOzKDJq699etmLDbB8pk/zj/D5NmhmcqpdJbhw1pK477K1eUwKm9K/JwEguPCoB
AI7cNrK0nnamBTp88P4tFh5n+cmiZtm9n4XccnfzGJOs9cmTWp2QrGe7uli23t4kEEJE/QdsUa5H
beiUkRwZswL9GGn/EhEhrRvi6Ifk5KQM7hTa5NpWKobKX+0ecV3B1dfp1Y71UUs5rBRpheTdrSsD
abp+2Sa3P8CKqzhKH4xSO/IN5sE+WpHi0IWtyd7EIxdWzCdI3hpgnNh2AejE2xx/brdVZHF/uGEr
nnal3M9WALTnRAIwbaVjBd+CfGirjWYjNn5l+dG8FZ0ClNun8d568GbyETlUs7Dx15+kIhCb7SZI
ElahJQR0IfepzzTAhpe+9F6edrr1veYXUTI1Vv6DprEAkHCVudx1DIOd57OlEl9owJGshVw63wjq
c9oeJalh4E9SBUgnahVyITAMR+1pCvHb/14WhRLP3J+atcF05XtuEKWe9PzZinbac9O+GyB+HvOh
YxIti7zKwkDKzwLnHm16ENMxDYnYu35C1309TKlNEgQVDrcZsksEkvwmhhvVhOyq4i+NdGotFCqF
jlr4DMxpFcZlnD9SHlOeFHVdOCGMH5jZrpn697iDSjXYKWdZldBgydJB/f6WZeA9LQiqwHDT9uM9
+F5HW8edd1H0nWcqCsEPT9SH9w54G4f75JZS3w85n0eFszMqDV7CzlHPG9brWs4xdxT2lBA9RZjv
8QieCdYwe5lCt3UI1/7wUWKSbiZvzNldNZYeYsVl386DMbSlYYhYwiyow1o8645iNRSGxLflvnlY
Ap1bULPNZEBZYQNxgvoL3RSAY8+hUlUxodaXOvrv+gOcelWQtdWyxPu/lXOU7XBwxoqQBuUkie27
BJSegBNbjQxCoLD+u71dpejN8FCNSmJahsCRkg+8+pqNy73LsnaCWbwUJmXBvcBWiiBacPbfuoMS
5/2dlx/cNJwhI5ATCJNFmaOAdyz6BcrEBfJx9GjJCf0xc+O9YFZ4s1bPf1tLPJ3Qlo2b18q2oMMf
UN2zqBtv45UjH+Zsvq3SdJPG6cPmv1FAYEA+yrvRd8V5zCSqnlN5uOKce2kOl0bLiBc3d4eqdzIJ
nXfWvUPVlMAH6SAzufTEJ+E8HF1vx+GoLoVheaFdcXPrhWMAy1rA9uBY9C5UCL0Y94pzqkPlD8Wo
p2kBcOCaDKr8iJIsRLS626OwX+NwTivZaZdA9xP9liGkj2w66ZWDKGZZsBRu2ElQOG/xMO+JawVt
8wBMctgKibmW4JJ6B3FuMkYrRQGT06TnmeiFp4enFY3T1xKP7BLiBu5N3E7LbnWcN5EEPbXZVFRK
dYempCYUWxFFNJibUV1Xa9R6Vbgwi0Me50/OcYPCot7xTWD9C5jX0hwlVxZ0KgqQrTJA75k4lYYe
7pu6O/e4sM9CJo9HPzv9DFScQ3e9qhAOFd7SyT/+u+xaTxnKoAYArDjj5R/+P/5RkzhOMS6Xv7S1
TQm9rNzqldFdIwwbb0VSqMt5f4g5fssEpG+T/YxyRX0QUvs2ZG6rG7WxKHSEOhcQ+Xrht/2yq2M9
6tfbm/ncpzkdLKRGZjUKuGWGZomvPiVBGIJFp6bsW5CPIgx81h6FVmX3jP5aH/F68d2ycDxzE+PT
IdlqHI6upIJfoVVJCYRfBULrPpwyNLQ0+eoC2vn0UodTfsWhrlKMD4HjYkovUO+25Va4gVPJiXAF
xQsaLF/+s1YZk4ZgtOKiUJoUPtof+L7eXlBuobbpxYQJl/E2W+BAHofxJLenDTUfAr25aVxnKCD5
xQMR/pr4LM0jotSrtRg39TV2msXTJV2vGcRwnfxQKTOGNiPl0hvkaK/OX//Ev/3r+WATuF571x/h
zWmw84BGBVCI7BgyGl7gMmBL27POTOkGyXXQh2giwh+kQI4lfS7C2Am1W1o7OKVEcl0bqZcviSk9
qp/RhghNx6iCBCY/ixXNZOyHKSJYCUv6b2wX8qL/MFufttQlywTo89SEbimRNa1OBHqxBCu4g8ac
J5weYeCbq2xKer4khfDcmbQF/3tK8UZonQ2bmfMWH4yLI/QHppZjBoCIM/2x9pGTgDsN5nL7MO2E
Mm/c7LNfDCGc20qv6it8f33DUlep4/vl5ek/5NAT4QQAW+EAVi1jeygz5uvALR/TBnnddbpOk77Q
M5QUlSY68icChVjS0RTe915pISxflvlzx5YagQWNF5w9SLJ6Rf+0RF+3SEgfQk51ZR7K6O1AauFV
w+TMau22YanSzf0qDw8Hu0CoIbgPwbJjtJq5KMdYouq+YkYCNz0ZGq1kav6p1NRK2PkLzUw/P4r6
ETjafmmCJBotipL0zoO6b0evTOGJ8tmBG7BOjhJbwOrdyRNytzQP76BR6xkU7CKxanBBuEHvgu9A
7KoZqbLEiC5z0Twqzn/J/d22BrtJxjwHZPOn+880UwENdebCPPRT855Z/UUdBEmJ5KnbDVa21kz9
tRyfPwPGUgTpPPZ2SUpSlzKgUOZ1WfO9OUoH04EvLQQy3SOq5iE9/vxMTXHMTanb8x+jLJzgOuNc
Z+aea4Gua+fklqAIUEUU5MK7Om9YTqCoguHrDsZ6mfyJZ8BqFIwqk1AtFfUYbn/0ESp6gG2jNPv7
RvBT/utT9R6lLVRfX8SqYMwx2OkMBeI4cCcGe21HfsYO5jGoZsIYzFp3RFRgLAxOU1RIG8hEYakg
mRITLiMEymdU1ikKjKx/Q21leF4gcbFQxIhwDwlu5W5Pt8aYRmK1ZGXvWiVnFZnf8OlGAGjZFXtu
MHQlozqdw/5S5JNn25nzKAZierFWdeRxixGafMjrQ6ZN0/o95B2SXRaGYBAKD4QSllG2IaFT6RWW
vr7pTeoO41Nqw4LzSHHBxn+CR3bkCjfBeHx0FQbTKAk7INTeoYg64Wmb0pjyvcX6rv+9jSnRm55c
KfZRy/8or03oNEQvZz2zCobXS7z75GdLpwFoF3tBdT6a3PlYTNdOHlieBtmeQ1e+2So4lJGwE9RK
+BXTgcYU8eNuoQv9XeGktpbuY6LCYc7qDDZL8E5dn2bjkMWULMyX/Z3mRCraUZphnU3SbgYV+aaJ
P1VcafaX869yhfQU6SKAK8Khngp1vUKHuqvjCxosfJLutQCcmfOX8ibn9uM/RfYJTi5f9SrBCZAY
mo1F+Vevik2D1dXIjLn5Ud70pLv2KL9V3cIGRX6jJ7hMLaNuvnF8sSo4jrhwktLqwFNJ8NrkjpKj
E/PhmGJu150XcniMmhOZNuBgwNFWtxRXRzpBAqXDcWuqOadIYrDSXd+yduzImll5wizwGwBxr61h
DUVz01WKiVMsFWudoPLkq7JZnQ4sK9ycZ2tn6FjROAWxsGj/s5etQFlNj+khov9+hUjzlgxNGPtS
jCpqYEgqy4sh1a/y1jT95oMbejba7jd+kiInslKJKfrYpIVMOCKvMCDl9rQQvYwjK5wWwmaoYxG7
SSxQw82BHOmQoVievoNxUPONGXLDIFx5nFnF8XYR7Zpq6atln5CQRoG8vh6/NjseEJ6Gznl0+z3I
eqbt067ljrbblB9LF5VeZl5s1zSOpxKtxLrfS28WCQ6ZgjLAmVKL01OZryIaFy9WJCTvxtHSRjdh
BL2obw6t06WHV/AfTOKXbIN0c9H+MjoxDQvjG/7UOQx1NukBMN/ZdH0X/2O4AaKZObQdru8AHbye
38OYR4OBWViebSSP/5PvrJZsJegy9+6iNE6ldAx8YpT7u7fm5HD/FMMxSd2jChpMfpN9QJ8MgdnF
+ElapbCinQZbQRhJ3VcMW2fMFtDNDrRMwNuU4AKnlv/lsbgIV//JsJw64AhFzs1sRIrPHei04szM
LPSikfBMs2jk0VER8qr6nly2u32HMdzwpFquSACEEK26fAOQrEzzNcgUGJerjX+T5rSL2UxHO5Rp
0wPKBGkld79VWd9MtNnTdg1uzaCBTvwOrW4Ll6zQEO+ncDm+4zUKBtGR23YW2Oh2iPDQhrs47Lq2
RMkd59tvo2GZ17P3Bvv0aO4S34etJsCOkL29e233c22hepWZ1WcW17kqPfDNGhnGS3CWWCqHuWJI
XoZ7LO9gZW3eoIogQI+aUlZ0InivvKnp0AEc7gIbHpt39su534EnIkPJPdbgagcAaL0UoPknK0vI
42SR/QzmVKHLqpHI09hmH6qW5Ty8PJhJ5Mlm+sT/PVj3SB3ymvfGHjuRaCJZtsmSJIi/ux0/rmJW
YauLpHfsXBhajwuS4VvW+NSD0pmhcOYD6jBODCVCFM9l8BJFnH/CBXdNgI7/oYsIsP9xMBOdB8L1
uMpt1NRqtUPOuuJ3X1kanPnTxpbaeADvEplN0PVe1vrDsQVw3lGptsgIn5qwHJcNW9zvC1UsMiWe
+7ylUSEBPI223aqfug0Rs6KH15o9LfsrquYiLE3UEgDvtFEal7Gd0961bJbMElSH3jq3eJnu1xJA
dQUyvEfpGhE4YOdGzo0F85U5BqWgRmY+l29LOW1UZwIv6LVJjBPmRZXDyi0G935Mq6FNO5lXNEZ4
fr1YyWvmJjKXO58rNWP2lYtQdLdwWR/nzpy5UVXAKdDLdN1HB1/aK0sarJvVRc0XTtCuGPNqvTOP
DOJDXd/rWPJ8DgYnDr2UbjL8IbC352LizuDsP9nXFNQYD6iT/2KZyKALRL/GXPuGLnBJ/tlHivVw
b/1GV7FknkQvN9j7lHVZCvz403L/M4xxgcG/mjMJZQbVM98tkoVEIzZuP8juVcurCcBGvyA9X9Zi
2X96EV/1eR+KyPD+OomInBjpF2evqKPOBLhH9dJJtz7f1ggpEvb5WE/QcZmMQ1GYu+1Y2phqBQe1
kcJHVgQkGIRlHTOwH7+xr1meA6nPq7WiJt3/mSVrWXICD0oMhlAvFw2olvmHhyjVKQ3ocs3F9Isr
2sXgeHqN2Ns6mJbqW7VkPMla5ysdLlGsAorcKZORAquVf9Ie7vbYgw08x62Mpz9pBqU67iW1EMK9
QwYsVOGHrhPxgb0rAmZXmA8uAJQiPPqtoGan1jJyhL7O9qYWEbUjiE30dqF4xACGFZAlQXqOelIf
zOZhQSTHHUte+qMxuQM3TfV9dNCsvQGe1iWxf2cgIewtspXZX7RJkBGlj5bvXYK/1NJPAig4h0Os
lT9gfCyiIf6h5V+nhkG382FXpNr8noGtBLYcjM2xPqh/1Y1iDQswEEOsxBhgFsNLCLUop8sRQ7lk
Hv4QRLSMMtyOU7iFZtyqDWX9Xho6rjQ+jg7L7YPrgP+KoH7BYvPUa2850E04mMOsxYgOsNAEFNOD
tT7bSc8vHpHeclrIi5+RAd7lyoH1dZSwOkXzCmGRI6yZ5F9FOVcwEsEhyKH3XRALso5YBcAXX+Xq
OmxzzgOI/7ACeqqrfv71273EwF6QA1QM0rlgFDEqKoGa9uCsn/tOmj7+qJ3L8vVDMG6fN4YRnOtx
ZnbOp69/NlLXNjXgoS4TmUtz8GoJpUdYg1SaJTEkulFXNDw8jEpBDOjHHuQBGHcJIw4jKd63RAId
FejkFBMHZJGNuzRNFQsyJ7BREy4b4wIOMV4tentZ6THbMpBXMhezQzCz5x2GV8LnMTXvcHz7inmy
OkQ5W81Nn+BXaIcDjePdUTxsrDlDVlnRdkginjO2HiEb+sPo5xiyofo/H7EGl6eH3tCj1K64OZBh
6Hs5dbpkHLXMxrCrbHcsSCTQswDg8LHm4Xpy17wqGII51C0Su3s5nP6cuOE3Wge63B9lySBwbfe5
yKgLZMtBOQR6Xrhd74lmvkDyhqe3x5TSwp5kHfH1s2GUgiuAZByHqhHePvriI9AbhE9Y0kGiyoCO
9P/brxVNk1PQWSqn0hNILmrfcYNFKx/ucHvhegkKkOK0AnaSzFZpodcNjDI9fGtqGztwX+StfE8q
BswTPGpOoEW64bRSAhwfAD2B5UEclGnGTLhptkfVI7MxFyIFgHH9CkFKuE8FGnHOZHW3yS90CPHX
JIgcnhvjd+Myu5yH68J+u/4CKgGKHxsUu2JrLHcdPskYVHMNx1LYoIZ70FeRg0s7Ex2T5aXVNvPk
1vSBIiB5cBk3lX61ZE96/k74OO5QcT5+tTCcSrdWTfBB7lzYuyzSxULXSeeoeyoD9z77n1mfr1zj
BggdovdDSZCgUoTbF1N6DseRUrSqsXjyxBRj8sf9MA13UFYGSCcLiO3bg83sfRdDaBvAR4s+mRFQ
WmSZyXcipbwdaTekNr5AIPWlmATVvuhLGNceLUKrI+6XxmkuJkp5ZAcunXJSbtEP80YQuzcmyCh1
womax4vODN/8HJP5rgSFhBVzP1u6nV5AoF50xA10ZJTjt/x/H7zKH8f+TRcXeaSpz6Yx/rlEJ7nX
HnC/85s7zZddPKN7Dz0kVyv6gbb5rFKXzDHOwrFC9G/uDo9ld0YUFR7+TYRySXQKf7fYLbLKoJLR
X/Tp5ymuB7KkUJyU8gvaKb+1jCpp29wNSn0llidG2vdh3bIk8DwNqiNeb6XkEAgav99HdRjCZtIi
q7di7IzWhVmVcZzgzDEa61pXi8h7E5louGHoMRlt8ifSkWdMo+WqklIeQh9eikUPjOc6vb47DTJD
78y63ovfBWX/ANE0BGTgI/wu/3qgjRjB5Fjo/uGFsN4bcmUz58xYKPEMtVD8RM2r1RXHqqUBwbTi
xhYIp6JJGx/46nwVWjYhWi0UsOHurAwwzSYJ5xeZmVGHvoOJabRGMOSsoZHsKZTUf+uTS/dCYfBI
BvXZo0gxwd+gr4XnePvC2AVcK6awPJjp5h0nFg+eKmP4oGhMtb8v5ZGydf8wGZfyqrnVQHNa6A24
veDF02P20GiVSM16HrFcF+2oH97HKfgDc+epjAGBbsblttPDSyZnFJaR+3I8yFQKuKzhRTdozEyJ
W0+5nLcAOwV4buPQHxm3u8gJ/ZWUI+lzsdYgtf8WUZ7iTuUjGLpQs4WCStEDLxi9Iuj3pmYRp2vI
uRYVlngEQDYn9S0GuLymCvAC6byPco0QadlW6pp4UBso9jn+80RhKjxq3tGKSksocRe3Le0Ju3DX
4Nj8AnevuUCkdri2uC00OHwKwBALtRFDLCbsidvgmKpKgSxkGj9Q0Ru0H4LGz2W9Nf5/iMt/xccC
Vmq9NnTs9C+tMIxqt5boHn4yMhxKZBkVIRfcCXhBsceiq5tKGSDWJoZz5ACei7oyIBH4JkTvMepu
99C3+aYS6K40GKXip1TPAFssCaBy5Eg+yzmVqwvyHRn/Totdq4hk/WoCBTZckxxhv6BGKWjWzjtf
ZqbE0KSywhLe2r+luBOiqWBky7nTDoVGPDQvghXK0gj4AzMyd6auEkUGRZw+IB+PKKQLr63MmQ9V
YI+xiPRlG0DByzKVwqHksYwOk9JAXNbPP5+r4kCPCf3zyAS0xDF1UDYDFyoF+HJgL2KE8VvZni4D
+zp9nTtlnk8ubySHXuAMi4pWpeBfXVNu4FeHH9adcVV2ywfceOeTWqTEWQwRZFbps1YbMlnf9QSo
ngFWpWyTfHtGnENr70N05hOQNwMTIa8RMHtgkqP41uExAmR72cQgsR8ROV9KkqIBj02R4kCwpDTk
ysY3+4BeL/GzdnKQ2z6SU7k4junJq6l5VQygelRZOvNZFsdgy6ocJKs0HTeKCkuRPlJbPMpztmGD
6MjMSV+m3tDtyHg+5PULBPoDWC+SlLiNuIIfJwiL98417rg4O78vgfiyfjI2b/e/Ao5H8HNtE4p9
5GWizjihcf9LumaDz0JpN7Xh7anG97GiB7BJM8OVEF4zP+Z78Q0TtwHz/CN3RCACIwwTDAysIw7r
R2uNq6Zd4XOqnxwwSAqiRf6aegyWeUJET8idkObFCP3p5PxtWYVOXhxqvYgNM0y3SYCH86BG7edb
BHq77gEkl34CertDJzrC1KDQnf7QjsO3e1UElULhqf2T3wFMuv7catiS8L7jF6xvQDPGF28uXt9w
0gf35ArRQUjbDsaYifIG0BFJAHQWeu2xOSNt553eZIep7pMzRnxfuSFBMUf1c0byWCjVi0QMITLA
FaP5gGE4A0Z/8tBVP8r48l7SRjtk0pHcxVOOc84wKLmuYVSDqRZkdjmK2BsBXgBLIE8IX5i5lEuZ
2YBzrhSqlbg/KsrkV3nnG+OMxa35jlqYYy608mjY/AHlpu2G0jEF6Rz+v4W74tEzDRCl42SWGSsE
S2eHuN9xKHagYl2sQ6vsozozbLDXXEwYPebY55TuRloUzlSx9MfK9zDh6R3xNlnzg8JT+2PMcVz3
q3KSZtGc9uhlt4lWJxpAyxGDKgXmlg02kXB9T7foWGPQtrJc/MkgEfP0tK+G0JtM+AAhuIwGOInC
ORjhfa+5E7rIbK0hJMc9r/gcg8Liwpx16h+jM2VJxit+XqpoUT5ePjT7LYuK8dASDgzHQ9Pv3MDe
ZOujvmny5aalgtGcAtDOF6wJnxaXnhuCFNYTOyKdRZqG8S6x1WMvcdOOXDKL5ptRgnEZaKQWwuyk
NxLubG4VFTC7jg63U8A2+RI4JvkGkBiOi9v9qxVgS9HCvdQ2T5WjNfahFwpd5PS1vK7KRH09HE2K
HftcTWm6LaoS3vo28fH2Yd/SFX3lCVb7uQXJrPvi24hgTTD1MXlRyfwvpmUEidW+SiivwdYRqyA4
J+7zed+NvQpGDcyY1SfMsBCGXoWGAMh11GoHzr7C5MP5S63Ye8Nm90XMLoAxUWIRKAR1PDfZwyLn
fUA0mtcmmMj0b6G7eS4Whv+VLZpViz0yTTY83yWsCUQdjQVeP0iz8hcvP1zfMbS30AMe2YBEiCjR
FOh4nXywDKhE0a0nksn9Kt4VGEg3/u8dhHjV47KViABJfVgJXkDRUCqr5ljlaRP6k6KfDtgibwTN
wS/AHxY4vy03dpa/TRaMj5GJNAjXAppioAbdUnsFwEfMo5J4KA7gZnotG/DHdUdQQ853BMKi6RYr
z3ZsveERaERndg4Dc4Qfj0nhzdf7xxjxy39SpsN25a2o7fcTGPWzl5rEyMmVMdSYWvXDSX6O7VQe
6n+6UQ7WxFji1l8nbHLiNOsAqC076b0Nwa3b5GCJmmFvndSzOTae1dHFJ9KQitts7z4Co47QVh8H
MfKeIRIw2qPGay3z7SnnH9vFKpUrgZeCKNUVqQxQTjwY5ZtWjFqF1q0WDm3nWhC7eqEL0oGFMg3c
Y5g6z7yGDgOMvZBSVE/dv53DpS0TF5cexZXx15guA1Jhwmo3d9LeZV/ZHuidi/0lvlzpAImuSrLn
S6DbiwgED0i0d8DUVsYN6iZ7S9nL9bYkb6k/HfFPoezqoRcd1ZNdodunhYa8O4hjJMShcyo5EjOE
aX29Ju203Tk0Y8Cz835GCXoC/MLYNMSYnqb3VZ0Hrmkwg1Sns62FF0qUL93TaU5HFJZ5P6lolZ/l
NmrCY2uWj95B8A6K3E6dTStdKGhS5/gvzuhsW+oqOLHe1uMoCq/nqYF2kgPJddmzhkT8jB2/So/h
uvXDIynqtacxzM5s8ag/ENrGPz/gV7t7Wu8SkszM7LT4xSPhWoTmqKqgRxSPFsydfV+7GKPtK5bI
zINmuQpKt0UU3YNfc5hLNQpwUzSYmoEa2rkFUGarVHDXm/M3hQvoWeQYM+4MDtgICjNsYDvxRwta
+Hq80V99hjQ/Yur+PCq+a8gzfyCJuAlJxdHsD37UZtKsSncgZKBk8XTdTwVB7t+GHNQOoGjLhR0X
tnAShVX2L+ScCx3VrMdRnf91p1yDoahhxjCbm2AWbUPs8YXGLhnou+im1ZnION6SGTA90SSlwhGu
yK5BRglRAPN3Qiyk0G7H4lVB3BEOTPQLSbPpN73E5LVgbvc6Vs8GRyZKgeiLGnmZ8G24g7jEKs1I
1p04xRdR2QXplPyOpljS0s1sNVuSLMa80J2t6BSFKxYMSTS0OpsoYFrKsJEN1O2QgZ52R800kIJr
q3sHyGn7CsbQHd8/Zvch47u/rm0xmQsbOC30BRdLHXynfGwX2dF3uQEhAAjkDoDYm3OR9J4cbWDT
PP4weCydT4YTKjYbiau7EdFDjs0JesaEYX8Uz2MikscVs6zHMg9zbEHBWMz1tQRQPCU3Vr04qUhF
ro1DaV6GHw0q1FhEeyd9SPYPLRCKJJc/rfC1zPNmGt9sDG9XwKgEAK/xgV7yKUplqQuSWcGPfG5q
SlSNQ/wr/YA1/f5srxUfwiNlzo3/yt48OKlmbKxSLNdCwLEukHrXIa+Xd/VlgqwUtoaNP+8YSwdk
zDYF/Y6x6tuaJJVd6/m5bQjojIfCbTeM8v+GFMkPpRbhVU/WD+aW+F8UdyTQ7zhW/eYvR17D3vDw
K1QpUdj+wQ70qy4t3ODd6Wiju71GmkI/CGKeqHaHDGQ7IqCb+sfi9HCzkIgc+PqeLDM32PO0/OiD
dTzj5RLpr3DS69EJxizbzcH35SHWlRQ61HQOzWmTyiS3vrAHt0CzJzdh5UYtyNOr06ACGG3gN0Pu
Gs4W+ZasPiwUI8t6LVu4S9tbTmrraL93EOLgFaFVkhwRiA9PVac4trFpjKhjvyj6cQw6xWecITdg
gy/beY2yz2g+UjdMopwNeGUH5UKaDDTr6i+69VDHZEts6b5McaF80oM04b7AymaX4KOI1MhedZf/
SrmbkyuPHo1w3Qg=
`protect end_protected
