-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
NktBronUy9z/j1uO5o5KjOqeH9ctIuiY4q/r4BKkZYgaCAo/bb/iCSawaT17/X9AqheJ7eyqkdHP
/vErcbvs7H+EJu3EP7D+DXO4ykk5Gm8hnOdrF1E6O+s04tyWFe9pGgeh53zWlRUkC6bV8sclvW33
ELEq09YDiKVTPcHxsoFIxA7fJEzyJpP8/nFdClAj7SeRzrmgay3GIxUQPN5vMN7M4Nw7VUZu/4SJ
tdnX38Eh+0RgruQuKO+zk1k+8452pmlKaBQ5bMM9kNbkczfjXYMQmvKvnGFGkdX6oOF+fikgnnZp
jpLZYHy5U7JuxyNDe8Jw49Nh9klhq0DUSNbTsQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3888)
`protect data_block
HNyrd78SLmBcN0htNSpsQ+WVb3JODqDY5NqvP86bzOq2u3Yiu6DiDpEoHb78KW1+HdG5jtklQo6r
1Rt1hLQwcQYERXC1ELVotkImErjGNO7R3pw+y9UOO4H0IRGkgQiss6uanm9hXAIfbxG1Ja8QjbuG
IeMk7ZfKUpspqGBrFmj+kcR6VZ0WlzQ+qNoroHCMMF/RfPBU7xLQHYAjWxVu+wm1y8BLZ0rtRWfu
nXPX9+FwuK4fPoHonjTNpcgjc+oBhsPKbbpQrcYS5JQO541GBwzTprleze5Dvw6k2YXbKjBJ/e+g
aDdox06A0JBpqWHrkb5nDq5rpNNz6p+IDL7cwOui+NdbYyyrL9b4k3XinlFSVaxklEB9/lsDQAuG
uXgtXRvt+sLCZuKenTfZe8OwGZ/QKNsGTl1CxxRt2l1p8RBsVeMNK7HMweIZKwF46n5SvC2fdMHv
5m+npVi+JTHk+4o6JwzecVD+hvELw6qMTk9B2vMy+S++P5XVU4qOd7cXgaUjoIpWp/PSmW1nyvza
SHPVj9zG3opx09qSmtMGMha3nOOcNaNLXr1sAYbMbWmKg0O9Et55PGcJPu9P/BytHs60TTKaSXtV
KMkvqNvaOuURQQfLQuCGxjTZyiPilUpNEEMXTtiJtcH93Sd6OUNCADrUTES6zUWuXeT5XajJhaEf
n1dN4NC/mo1YzwT5JMdWD3PD8ToexR/0Q5/Zhf9lVbii6vg7MDXoANzUEqcZ5EPhGl9UdQvcdKh6
jUy1BZHUV6fiOMvab4wBAA6ORzXCpMGxrAk57R0NysCieQKTq2N4tuYil++3De1OVjrJN0s0Lg09
xrGU0v2NAVDedSj87PAlxl+j7vuiDM72dcuuJm1zIK9e2uq7Y4jAbLrpjdPTBJ4KU8aTAwkKQt5J
6jV504snLnSt78JU660gEwMKgZc8Tt60Bh1TttbcQ/KeYlFw4tpfPzhbJx+1p6pPWYwvkHQ8zqsN
o5tT4XN2CxUEJzqPLuXyAvFwcCsQ30W3BB+S1SyFYEAn+ZPHUqpxMYEreMp2fNQULuKoEQE6/YyJ
thCmJyjZ73Kp3RFpwk3arnp7+s7fwElLUv5HZjSpX/NHb4zV4hfdc9gODBtRsAVPsyzXt+VJWpqS
R5V5ofr6ceh3mYcRysvz9MFc/cABihrncnpre5BbnvpMmq0KuBuPA0xm+WUT5vhmt+K+AChcqCaM
HX2GU5EdCiJZCvBHiLqI9pr3IH5hYrraaHKqNOLL+FOu+naVwWCI09FVZuiZnq/QZnHEMPCHB0Fe
w/LdBn2KCPUBMsgs94x2zPuKiBKfdMdkSbBBQy2fecq0BhD8SCA0O51zTROPoxda5TTEGC2VZOzU
GPNFV2WmN7QtHssbA1gM7lFQru0b9AWS9RzeqigIJa54FRK9V6KUxTKbvKf0e+3jCsBmitp10lEM
R7s4kKcpSzTZyOSZPLXFCp7Uy2xsRIeCC3VznK67a5K8Uh9HQP9yBmMyCM4huoCyL6KXfdtAdP0b
YAwga3RVQW5Yqtz0i/32pK46keHsrQMFfEbZDq5zal+r9DdTrnSjzThTzk8Wbwc3w2uMTaS45rQp
sJ3Sn9sI7HK1YNyNp0/gsvxeQFxsrUlgf199Ilhbi9Mcs2XfwefrmCnN1/pDzkau02bJYjSpi+P5
A/rrUAadITwOBHahvKO09E30azRfD3sIohSZPYkI9Z+PkAep4/8WvYbBjQ7B4dpr5T9bwmKry9Cn
d6+nq7k9kPW1JNQvDFPZrJj5TCE4U6aTwyh6iifYQIbGdp/veRaT5vwtrcE8CRgCia9lapOXEBjW
/1coQc3IdhnYkEbT8W2Reefjs0Umso2eDByS9WwwC4qwaZqJiRmmDkT3flTIVhZYQFSUynRkuU8n
/pVOcO9ZJj6fWjXX0dMyn1dlx0ORZWtEdYzKRoGdMT7kIy4gEJjGBYC30y2gmlPgA0lsPcPUK/ab
3U51nkdTot3TYA6jo4Vr1MuSOXcbES2GSkq3nfRLFNw6UQ4G+p0yJV0DMHetjPo+e6XQUYTnqHUM
PDG9zjMnXJjH5pYBG61APD28+r3Yo6DI0kYnNZtEf8v6CvmzyyXPMIcS63u3A2p0G1LxzQ/0xMbM
qpP43pKUDQlg7ixRdAzjBSv+TNVk0m3yO8yMlXKOIuWk8czZqeOasPaYR4NP8InSJPP02pnttex8
2C7IvQdZCM+clBqMHXJC5nZHCZaHWswd6deIHpN6v91/f+lhzg5/ZUVwX9yBWd/BlODlMdQ80HAL
PuZzLmqubyFk3wyvC/6D0HPHwa+ugVRJxkeUCNw4jlIeAwLHW89AcZOx6V6YmS7UXLKSY68n2d2U
UyRbbg7FTEaMF4ugbaOb7IaMOtHuuTlvs+R2eJe9O79Rxgjl5r+IiiobqBTPqzdb2oPhlQ1Pl7Py
RC5b2ruh5/eZYpTzXhiXI4hiRNJ9OjZY4L98tn8BhFNKKltu8PTnF1FQ/E7XB4IWu++JobyUo6tt
p/xYiwzQqqmmkXF3gWGDLLcvXMywQGv5TrHkTywCh5XGV/dcpy2OLt1LWLzRzXqt8+ztEnljmt9j
3EHlxNdck0pgkjveDyKevfdo8mEUr86JJc/bDTiB+nOsMbg1gsK33+NZjfN19Xs7iujJ76xKJVeS
lUhas5X3+BWPaIL1GlT2X0tKkGAZIKCVSPvfEPE77aJt35/YL4iOQojTyNm2S3ZV19v6D+FofYma
tRq0LrCIOt8AzBGouNwF0ADhrSKxzyNbhlLRCLTcH/w8fHkUXW7ZNJr/nYF4Q2XOAWsiTzhJIXTn
VTs9TTEjpoTcd09PmZ44q8cGUjNAJxKxxmAhePgkQ05r6Te//fhegXor/Sf722MZ3bEBSmf+0mRm
sx/a1hz0v7cVOu6OOzUDWIt0o5iqMFM7oSe0+/YvhxAzhi7tEWPcXgGw2M97uzHu13a91aPCyiE3
E9wm6ve32uX1/5mZN6QcRfawzClVKbtuwsng5rKRHjqEXGRksBx7pzT6wNITyqLFma7O2T1eF/Cx
fsmK9c1if+VzKXx7MKF/WEo8rayMJHqUP4vFLtNDQeqn/kpMXpc1pe33mqXIyev/SIaefWUrwZC3
CLstwzwzx2ip6SipSBv3wtODLhZMQGf/7/iWDc/FODHZVrLIak9oNPKzf1M3fgvbpA52oJYCGK2A
7tjb8Pt39OUucDgFxELHX9cCpjbNY8pl2t0mD3hhZk9vInBITeisEVhtENq8nTUdt9+1r0mvkJRp
H+RRBYSFtmMMIlFp9sShKGPwhcx/9LYddV5ZzOt5Bdzsbyw42yfd2TrAk0YmXUidXhYmoy060UUa
O62TT88RWB1Vnssh2uasWAMfg909sFcxhlunjEoFUCTXIrp4caj0cNM/b72TOwQXupP4fp9B4gSY
sGdgizgcz2ZlQw586v0sn+6nvbjLLL8o55HYQv5c+c39wndK8ikpTvDEQUVMgbTHdAGOLLi4N5/C
n5supnBSnro5bo6VC2Fg6flq3KN8rE7F+1cnWtKr8zniaT4YCv8p02K1DDuQgzVzInVRayNxi11t
GsJcUN1hZ/ZSMHgYKSJ0jnGZlri8fD8G8WMLiXSaHyVsgoWvU9WPfTtYc1bISvEYGdQulXtVvgRd
pMryvcSrZaofMoJAqv+prPc/b+bXVOlurXNT4KNFBcpJhZ79jpgF0YFw8NIlx+ZUC+teOJM6BpBe
Zo0faY1V35X/XRVizBiw03YD9AyAuvR8Bq422pfTAv2E54pnSGb8d00Fa+bmCdgq17ytOPcg2Fsh
KiS0pyogOSih6O31Mg+ZTmn8xHpl9CRZ7H+jD4Ta70g0iNp+hiYrpnhCRdvtAVx42H6QOgYagreJ
lnHSM4Bqhx29OsQYhZODhQH4QmfdJvRhZ9BclOLXgbV/Tzuf/+geUy66IxOeYrhQ0CM8xzNqlsHD
DmZRBirhe7qrIQZ7AnGIkgUM7Ecj3+SwlQyFY5clLE+4q9bp8aZoH63wkQqPhFb7XN0ZsGMbQSIt
ZzqogFN5ppu7EOig/lyzWL2fez9fHe+jc7TY35tP4SPOdfwg+blOFGIQbMazujLD0h5tvZ49MSDZ
WKqMSnYSwY/w89Ers4CyRrGYXG3i5+/TkgmFe86uU7gRxwOAony5MXf3qpYo607oDN521fZ6+OHk
IBaG/lAHJAd5KI8nkbH9QGvnmZFmFeIfqENyKR31feAGb530leg+JvkUJLcmBhEkmq0GOSVGUNvj
L5BPpjsBxzmdeSK8IodDbAoKaRcvfOmnYDDGgPAiw8EHI+RFtWnNL5Wk3TAh0MipdErxFdz9PzxS
QMttH4MyXu4crbcelJkbgIXQ6de2bRZtxGUixT+Qr60vN7KRk/QiqkcD+giKgYstrRAxYxXqsJQx
lFWTNj8jopO31oyX+FhJVj1I75vARcmVWtRXgVl00XJ3DksONt1V03dpl0gG9qEeEeFPk9A7FmH/
nslvE+3uaMGNxW6FsJBm/GI11XkjW64jZhIyBoQRei0Q97+VP5VudyiPXPCzI842M/htDKVwoikH
p6dwacc2MeoFYoQVES05pgGbfVmcVgegLB0rSat/rUI+R85ueu8YYaT2F+L7k14RTuH52lO2951R
/oWYC9Wa5Cv7351mER3wb4X18877McsyF6LrPhIdeL8HZGDLhscTFLvo9XYEGBB4gzXi/6ogG7BV
ojSIG8fiLQ6D8JnBcMUoAxBzAmi3/Tpbt7dT838aZPzFgC0orwt4TJvdr7UjQtGWZTIkSM/TTxqs
dLautRCizfZ1WJKiGwZuEbm1pi+mEmaAEveThNySrEgiWE75ufSQmzEihyn9MFiscn7y4ObV2YSN
/QhakZ6JOYSZw+b4QmltDFwtkKhfslmftWlr5a2gI7K8p6Xa/smi7pvUiwkbbID2r2oPzdYcCgPX
sjcdCJ+Qx+vYv/Nl3WralPjAquDosxhq5Zu1yxb2i125VLkjik5/EkBoyPtLKXWByVAVznut65Wj
S0FJFpUItW3xiuTM70auSpF2aq41Tc04RZByCFc2KmoAkuT8qeREDqYjoqAYa7bHEQXgZkQ1igLq
xassBuySl9cE3DgSXI6T3z0jSfuzbHhm4qSY8nFIeHxlsKL5Y5xA728dQ47Mln7ZNlEbYTttMcAt
63fQgdcaxR+w8hiU
`protect end_protected
