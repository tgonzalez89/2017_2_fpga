��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR���[{�T���CK��TC,���:�
&��d!��]9�'D`�"9 S%�aQ�`!�6������V�W�l�a锦E(�\gC�slu�4U5=1�N�m��l�9ў��P���B�@+yg+H����Q�����v�Y:���NS�%S��S�@,�^���Y9  ��^�˙��F��3U����`�j0S��O!�,�g�)׃=�`(�h�'{��E~pVʣ�j�)P�J����$4ަ��ܓ�p�V՛���Pu£����![��S�퉞��\�� g�x�> S�
�hN�('�'��]4g]�$�'.�k@N�oY��!��L�0���3U+ ^�.�0� �r()ן��6�m��~g�i[u��}���B��?�E;����*�E����T���Y ��a�׼๣|�"���.$���e����X{�&��u��Ԍ28�z��4�V�4Z�7f*��$�J�yf\��)`B��3fE�SR�#`��lޔ�����{+K8l�����r`��g�b�s�Jp~A���==H�9hK�>��Ka[�t�Gʵ9��<7]�ܐv�UV�5r�������R;�(j<eIT4�p�e�S��	k�!!4�L����W$�T�����E �)�e��E�y��/U'���H��1*�l��f��e���Z��%����֭;o`γ���n�F찕�^��5DR�q=5��KR
��̣���E!�Fz��tzb�RO�s�4�W#��N�I�Eݔ����h��j�)�5A��K��Wz�D.�3o�?��J�PJ_+'PN�V�.�3�ڻV1#�t����)��`ʧ��秏k�e�{����iwEZ�\J)�}܆�:-N�ah�h���=�DS/��F2B]��
�s���Σ79f��J �c�/��Z=��d���O@��i��G��	}gn	>쁏��4 �%���+V��b��a$�k��+��!��V��F`����:s 8;4��K����_G�Q��/���'D�)z�d���B��˚s�*���@�_!��xQ�x5<�
b���s��G`�IU۔���}�q�ʐY��ެ&��CĪ~#|�&�i�i����%�̘#����~bC��5�*>�T�E f�^��������u�l�� ��Bf�%,\���(Qf���� նL^��"YQt�[�=��V��t�ԧ#2�*_��A�kT"��"g�<t[�|v��|���_L��_2u1�p�w�;��uhV.�ٙ����`������hULM�$�(t���SK���,��#<(*G�ށ���[�����j�uB߆��I.���]U�z�'�Q������nq]���M�:E3wT�L��wPKtb������sD���J�V8���^=��,yB�v�������1G���ͭ�!�q�{X^�����华j��b �|&/�����(^�OC�y���)�1���[Cw r�"��\0|C�f����>�Eב("*��Nx|r	6�S@H�kq����5��h�r�b�O����4Ş�Q�r�5���Q	�^i�c�0�49.g7�e)��4j�g�v��~O��N���c��7��D�`���5�-�b�NG������WbrzqJ�.Lg��_L�>��_ӑ�������
� kz���-Y�(�{\�F��^e<���&:��F� 
�!l�#r���%+g��S���o���1@����#�4��|���.96ͅ�3�Zwl"5h�'\p~����[p�@��Ԉ�*c��v�������}�"g^���;��7b�8���(�ӹ�iL�,�[ �É>S�A��9�Dؠ�ӉC$�8�_Ы��z�)o���ʗ�T���NrMw���ew�=�Dǋݨ�z)�ETr���A��E��"P ���睤V���e�O�28!2���t�8�w�SE:���~��r"��V�38���z�xQ�ګN�qi���W��m=$��e@tܞ�o������F��q���U��Z�u�R�lOC���%׃u��s��,�W7ZS<h:�=!�q�R����Q�ѧ��!c_d��r�TJ+��Û����q��Ѹտ�"���ODDC���F�0�|n(b��,�FA�V�Vn�6@�(����i�U�K5�)��v\�k(}�܅�Me���Bޫ������(2�3^)y�;���K'W�Et-�G��YH~ﭚoO5�ְܗU�fc��6嘥�\l��5ۑ��:8#���u�SǓ�yH�*���Y����
y�g������8^�	ߠ�_��v�0t�!F�-���