��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,�Q����ф�74$~�I#���F��e�.�j�7E7:?��6ۘ�:*&	�ipc���b#%��	�A�� ��0��'g�-�ṱ�3q�V�ڦ�������� �W^�U�|�B��|��w�rNu�vZ[ZwŤ�i�2�3B�!����b��c�c�[�e�4}�T���p�.�2(����o�^0tu,%��g��s3�,�f�UK�I�"�G��`m_�Y&xZv�a�����R{��l���똠d;����׭i���.�v���y��6�Â�@˞�N���$!�i����x�⹐t�ɘ�㙚�b�/0�7������d�%�ڀ��d�%���	{��~h��TP�t� Y��SK��5�;��§���ݕ4�?�r7!q��d^=]�>C�٠@E��B��ZO�%��'�d����*�B��,��	(�>c���]�l@����6�I�?t��f�G��bև6���"\S�{���e�8��U��$��к���2)�(]4�X;й���Z#�;��&&%,e'���:TM�D��������K���Mн_Xÿ�[d[3�v�rN�l�x���nbp�e
�r�4��'� ����Bm�ڛUz|ԅ�/%i�l��vySN��x�,��u���Y�'�J�sZ~-�Y�OM��Â��XI`@7K�z]��OH��5S?��xd�] �頻>�����\vI��?,�j�鋊E/�v�JD�:U�Kj�P0��s�]�5�5��7�^C	���	�cUh���$d� zn��30����t
:uN�=��y��'�|]n�Ti�fzA��Ɩ�x!^�}`��+^�	Iv`@͚��$O��l"�~j]��$�'	���ѓ��r�W�7^ڰh7���Ow:�Ȃ� o��TfwE�I3�X3���R3���g_1{N�Zs�?��z�]%k?|��:�b(KP]J}�8����b����m�)�|�Q3^���b#�V����	�qב�Lbr�M�
~�-�|���S�=�����E���h7<�u,c�D=�Ρ)A�,e��-<�ͼ=��>F\q�$d5�Y�L)�#dS��3�W�k ��!!��C$���C��`J�~�;E�x!z�T�c�����kVb��0��'Tt�Ϊ�H^9�;�m�eJN��Y9^is)C��Ǚ'�Z�?�Q��t�R",-��qUP89	���	���t�����Ӏ�>z#.����q���&� ����ܰ�h3�?a��3k�b��O�5��7Ĩ,�O�x�޲����4��\abv����?[Z����~��k�#�<��m�[��I��#��d^��E@<]_�f,~�ӐBߋ�gF�R�_����e�b�T�����`�ĭ*]-w���F���i�<<��]~F�i�u�|� 7w�"�a!��=o���U ��t@/VYC�\Z��N�.gļ��4�������t�d��_*��Q�5��Zj�v+��*f��ٗ~J�< ��;+w���N*��wD �,��n;�-����V��M�A*x2�4��o�+%a�D
:��@������Nf�T���e�����HQs�z����q 】�5��ܽ]�7�7qC�Ɔ4'�C��/�0n���E��$��V.x4Y�����IN��?���hQ$}i$��q��K:�{^6���B�\Ϸ��h�%p�"��C��L���+����� pXnǍv��ao��Q�	���]�����
�������X�л\ϓf��ٛo3`�B�a,�\�_�l9�>[��5�b�^����8��G^4?�?�&O�Z�eo�5eiN�tBs���=�h�~�1UqY���	�6I�r{�5������`}�,��i=�S-��dJƂ�@� KQ�c}�����0s�y��\ݻ0��JGV6Y���ע �L�D��O:M�Z���^M�y�2�2��S5�_�XU��كE���\��c"�=��x�C�Xk������A�ش0\��>�arpQ���j�¤6�ps��:����Eﲹ�ȃ�H��h�X����4�V�l�@)��m�:��S��&�����h���}pdo9��v�#NAY	�^ئ�\��a��R�;>e��D�l�A>~z	���