-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
FW2klCr9BAUgUOwOED4TpaxAvyZ1xMIk8ZfIZs9zXr10b1r3PlFO1aOG/bCydhqVEOz+6NnGfpxN
aHdjwy/JFi1TNCzW1AMFKSXLUxg9sJVnVTYp9lRTMscYdEZ9ywcWsFVwjBvPQqVXsiIbNzzRJObO
+/UvPIUlCFPIlxHnRzyQs5Mnf2tH8YIUXS5Ll28dYPxn6A0U0/pRm3916hzYrqgz5wBE+mGN3+P+
col38g574c2dFxgOXyxFqaRnTUIhWeqKQm5VzpbycK2VsYLVHL0pRJZh9QjCtd3zUc1aKwrdkeC0
vktcwwsT244OhFemB6XDiNVyq1Ng1hUHS+i1LA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 25312)
`protect data_block
HZ4cDdFmTqhi42bT9x0QVpi1fWVH7O2t0Gb+/qz+DQPa42I+inQPsPUjBFKw+jtejY0npboMZVil
QiTXjVwyd27VOFRcl3pq1X3wyc/w+MlBS8FqGl1GreCxRXNDPZ+FGbYEa8iZmIIu2Zx7sosSbF9l
Jfwhc98JpinFcuWruV8o2lSnnv/UilEAGAx7JjcgWtWKWmjnOPSVJGW3Zawb979xpFr+FXhXYjMl
p/LfodIIapQrEB3hCD0ajLuHW33At9Es/PMn2fzPJNL2jE2kW2hPZLRFcoFO1PVcbukwr3fso4A3
3MP73WliuSbpKD8JzhxmZPE97dYqEyIjtdULor8pJB1yf9EKIDXghSgo3lPRUu28SO8BwHz4XQRr
mZd3tRBc68bj73yrf6/6Zv68dVz9YUp4uQ1AxERp4L0ajXCsrlG6bfhiyF7asp80kQ8M+Oiw8Trf
ffoGJjaCwZ2eQ0uDEgLFgL5ngM1W69YmPI7+pmgox5+DUnvzBpaS5AtiJORgePp1cimka86l+ZlO
Y9zLBA11JK+vkCLitwS4RbWmm59uWeoChbTGUmqbnOCWtEuIfhhG1OG9JHS0VV8uHwCla3lX+Fvo
p3J0pbLCFZMkfbn0JZFaNbFDu6gllm8mah/CXSL00Hy0KYnXomu5RKOEJgmD4rERVHLQ273lNGy9
BO4rNtnARjBhO5RwFEiivTINvQxdZiQBDqTgSCEaXfqhJEBfD0VG9vSKVHl+kcp8twsi01kTwRX9
NMdPZKX+3eIJHhRh/hT7J47/7mtEH0Z5x42KiMhLYXxGUH1dNfDHrr1Mgvnj7TRuJUnEQSpWzMEb
g+TTnEc9vWGnFmV6aqjDyyaaqHZQUXfaGdirOE2hb7t7PCxbpbWaDBA/5NblFeJUcaJjGpaTt2Zz
8gfyfVsXOiYTZJT9pAWlYmz8BPaIIGB5Jz/c2D+8imcvfKN+i4qO8GaYo/M4Ny8bs1INfzgXfEWT
On/UbPpr3SnN5gcQludf5ZsvdkZiVzqRBDn9Ye5Zvi55qDzP8PcMctwEDq3eIpfggHMsSSIB/jud
Whlq369SdTO1+PL9g2HZG4BSjkAQN4wVgcTmBT6ruEpgRq6mJwnhT5o4TiiN0OOmhsbTI31wytNf
GUts3eFyvYg8z8cr4EEwdY0T3BAqu4WO6D6xfN9MZ0lgBu0lTQjQgbYrUV6lQW3Cw9ECGRlzw9lQ
zsUdsiGj1kxx3n3OwP8YOHQNOitW3t+YPrt/4cY2kNiqeGgI288UMVg7e0yx0+7BVcEH6Q92Xydd
3haBhEDEDQABJGkffqlF0PAA4c+hnJOfyCE0w4cxqMOreK4+Fr0AAD6r/yghrYgzRDkajqmvTE2Y
/6d8wzhezuqNCcZBOTsjlNX6LbMTRBjuJBG053/jET3w5gbDWa1bl/ttX10f/f4Oc40T6Jipemw4
vDpkMZhHeuDsxyGTwvyFDv5BJnLeqRCgeiJ+sqEQZv96hltOmuopiVtuKwV4rLWGk4tmTGKmHX2E
pv6lDQsBTW7ovsbH2pyyB64xg87HlI6Lk5q/oCABhVAX2zGTBK88LHHKIJHjnsASI4xBlPnPkfbN
6SnbmmaRDCcsv/jPLGndcCV1yWMJBp2JpATmpG/eAJApcAI2WmZm9bPtrhQ6OM7R4DVg2NWN9S/Z
yuuIVpTzmRnx/624AL/f4Yqcju1cQlZ630YA3YuSGbXRPlrql5F996Ianyt5uZyFr377UrkhFWtt
bosBnq7TdoggFrH74Radb8g8ttYkPB6XDSIPijpERv1tMlkDD8wuzLYKkvtMTRAqHdR1s2RNteiW
wfY3uH0/A889RQ6gElWYWjbsjv9T5amS82Qduzz9kq2IaP2rYKqDbmKMiWV114qiv0YdAsdTJUHv
ucnk6tRQwR8h40zLp+j4oe3p1JkFgtpQyXAjZu1T1tf22hOqjE94q9joHPtzRJe269SltD5h0w3F
Ep/7NIreKPJdmETK8/J6kgl3wP1lDTirqWVNCJk/ePR4j+93WoJtMFoBxVGMrcsNuwCPGEd/IW3u
/0Bv2hVRN96lGSDtajeArghgDeFdW9CLY0tvFXy9SnDxmcmYKiwRuJMYzs8BpGrYfAEfrNsEKPuR
bA6q/axACCAuudI9aOlb7Cf5o7t/gurvcC0Sc71MaBVnI7qVk3iMzQynwbh6GMItFp1yUj3JAIAM
Eyg9MOarlThiwO0Z3zxeAQooIwpJMC+1j7rxM2602HFkinU2cEkXnnP1X+HLCCqlsRyIi4Uwofza
ajBfO358aw2Vd9TLwlRJuyx69YssA8dS1995thT/SlzRPENLUBW1JSxnCQb47iMKVJBRg9Du9N9w
AF6lCyVG5rrok78vRZpmvu/BHX4Va7jHDTPeiaqh6GPTtPNU8hHDPG3bzeMcytgiPmH+xvFTmjax
A6TUvffVZNjeHpPD22nQvXPjjHYYHsnFkRXj010wk4YUvR/+LaJcZsrnoJhOEuk8VCuhaaxvV3vS
DihQqG4HrXuFGLOiTIrrax93WkFuR0jDGZwYcQtwKUSujw1Du/Esl9bs8cZAu17y1sdgP0rheEcN
PvLNrKR7lPgM+zT2sz2iAyIgWfleJ58Fj9flAX+jChU+xYMgam5LaU1DjiUtvL9uvrO3WxPdSfyJ
9GIGpcQKStYlC5XN2Urp8GYR7ubQsa9R9Ec5BP+gmWneLX0KbGULdcmYXpFrizMNHBCU05i7EJ9G
+D+5so0LefLbIKcPsySpCQN00/2DpJY03DvXGPUymDT7t2sFvN2tvfia5fTAaMGQXe3b/LnUjrfZ
wiX2rEM0/i8kD4o28q3HnhVdmf0/5qCHQKXFYiFN2CGZyNqPkn3ySiWxtsLD6Q9EXRPBQ3pSTnWx
5+Kb22crse6ddP6i6miTmPyB4AYg3FVpKUvHPDgHkeiHZbTvI0bn/Wv2cft6BxatBQ1VwL72GkyL
7GTYAwzKuUAKMzqPw0k3OXMpp4ooREgTWvnNKRwq/coKDdRW93arNnA5M1KamnmNSugGkdQCev9J
W7+Qq9lPjtTk+DsjtvxsWvbCMBUOf41xmPterdZdH3sEap1JSI1OmAx+1aOHErOpS1R3JDnmgCOG
eJjhjkhowabQ0KjW2JUrThwO5eY3Wl2v+6W7rI7JaD00LIA6SDM3hoJ8f2unj0uI0PJ/UwU6xpyD
bhhEHQHOZ+JnnkuQ+RSWudAr2B2o7RNZN5cnZW/RgNgfHU/lw0Jq5rJVp87UZQcOyeMv0ujvzaNZ
3G2STn9S02osO//+g675vhbTVOrf0xMfdyWa95T8MuBS3d4sEDpdZ93qk+qSjTGpK6FpSFqZePO4
cWVxML3ZXTn92QRwxzxoe9Qi14zJTBWZKgWuA8F0ArKVISIgGTVvbdEcQ/tU8noUIhLsY3RqEec+
fb4BFD438p6bhf45kDDz3w4cSax55fd2aOe9MavrhiAY+sAMSOi5QDThFGo6Zl2mvgo+TT/Xyf68
zLNpWbAunvQ5DFg66hJjEjXAKiC9GCnbGLIt53FtmBRUKZutrPpF3L9rdTw8kUKw8q5cCl2t7Ntn
8gYTxovAELvV3hzUbC04LAEYf9dUz8/nOTSqi3xWnkS0O7LnXxg/sgeJVATWdk8oqDcMk5OtNwBN
27KPn0Ae/IAtAqNhtlpKA3RoIw5MHQzQUU0GjrPTZfUI//DcMy5a/gXXK5JcFPFWZS+Jo1agrtKJ
ahECvDaMxuYvw0M/oXFWESdxrNPm78AQxZzeI1URTVc4QF9Kd3Slch0KtzAs3RG3SwC7ItdmRoYk
F/rgLc1krjvgUJkDouQ5H/Rf75/1O6mGxfsBmSztitsSXZrYKxqyJc0JWK4olw5Lb0qDb+pR0uRX
zmVLKS8IGdHjCzLthyt31awD7+2fYLs6wjVXFUw42qvdU/PtcTygLS6YNqdyTxLVpmuJ53oOBaJ/
AR9k2nOa92ADL3IeNM7jzrKL1q838qcJUU2Zr27t9iClM78t2sK9PlKEx4/d1tVe7oHorq70z7GD
ujPBGYPoEtmIIsw5am1RsQZoMSMkWEDSUhzoBSP1bKrVrA284ju+Eeu7rIMX9R2tYutvqmnAxdie
thLDKo9/IaDgcvR1g2ckAkGv0bApl3DB5OpCMrr96T6r1vW/vjHomuiL6DrscrbuOoTkp1JVTwWj
7xiO9n03DNB8yF/ag1cbJbQl9r5i8VrHwM6/XkiZimVOvIsXIcW/FSrLEfqIfDz6pb0CR9hCxY2E
4o0KelQQ92pfPha8dlqjeTaOAe0ktMkC9ROME2gY1XeYbXAcio3DBeFbuAyMiF7d1nN00iKk0s/+
y/oAsUxnPLuU9eIpUkPTrE/sYwVr6pB+h4kaTgF6CLJbtdlcACCIJUYdLtOFMYBOFEPiijquCokE
2IX5R/RuupwAirIg7ZTwGeqEGQSAHRLLqIHeEaUj5Eo44kXFemNukpnPQMeR3W+Wwnu7RcE6GKkL
r4Qf14lOZ8cr5165S6F1CbBTISOIsNJ5yebyVKQ5O+gDVCU1a6kv5fmBW55CtDZyGLNBhYcjkigB
2t+BCWuyXAIn5vRq8/clLESGhg7JIsLJ8vhPonA8DZF2Qox9gzbxH+fvgBMJadapM1B8Jz2ksm/L
CoHdxRTTHC1Hz7gKH2vNhcwnHneMybpeZyvMSezlu/4SkEldqkQcNS5QMyAnIwkEq9w3Fs2qPz5k
crzj35o40cKfvVGby11dSSrFw3LvtRXrxMpN8yrOIfCOeoD3zURMWVVot4VeJpESxtEvf7WIY/Tr
Ktj29XvqiwNffy/k26d0ef9gSfR1sYxgf7yJBp3tQLqElZwf3g0iALA9KV/yVtBvk045nCDbgqBt
HGysgPXsJhycAF/4Yg+dPs5JXeNWKr58BC/OtwPxKaaHxZtAkK6ZYL5gtyNefhZEI7uF7VUccLKR
yUMNdRcZ2fM8vUl648kvOyEjVL6D29kUkqCnZ1HfwSwqmFJW+BW3g2YC+JwUuWCvBnrnn5SOoacv
sdQ7XuRUc1A8F7Z1m8dHuDxVzP+TtF6ZyVmy3J0gXmSarub5/9B3LraGe0ODXZclspA9iD+m9UOq
ls8swHxrYSNWFQK6xLFjjZmtZAzCy7PX1A24hSycYgG2LvPmies/o+RTa8r2dBKjSSkrlNqVGSsC
2tge8iD+3Piey43fVYMh8byk6/9MOkzquTxAl3j4Sg941pNmtX6ZQSaBGdMUBJMUhRfqtB2S26rl
O1nvYzFoD/KKZsY5chSGPorVB7RbcYtzfB1sBpM4PMiwYAjD/2Ka+gZl0rTOubnSjZPZxjd504/k
gUBJfBz/XcDDKgBjPApbT5y5RRmL/ukKQeS1AR0tbRyJ7glCogonxV/FnnfV1vXRKgmfXBCyHn8G
cm3B/rIZSS3X5GYOHkk/WUcJhxM13/t2W5MLLCQ3GPIOytopzhG9V4SlJ2fnY7ITgJ7I3u+4ullF
JyoJ9mfgrETuk0xQC18H8i8ExNh1ZogYfx50CdYn0RxGMNxkTUu2GZTVdJpf9Icmcmv9KZHnyWg9
mrSm5ck33H6zH5bwy+QYAxAZMtnhnO5OYLByo9q0XtuNZGt5wQAghOxbaM2rHpZK3lSijP0iIoy1
N3+EDu/Tx6wksJbL/3Le2RN4Sl7ARP452psGwzizHBN84ovnAhDcnnv8tDNBCcoAxztYiHe3tkIs
VdzwSsy8B1JtLVO2gMsttgV5uAOyJJ0Eg+3bWC/hO+ZyAHCCTtkhS3M8mrN1CEVU+KbGzafiYtrB
RJJ6y6lhqxrrx95tKRRYa1qpLFLNZXkI8td1vHbAwdsACyn2rrOGPlwHuBIzbrV72j/N2VM1x4/B
V3jrIBxBYkr5SfPI078Ete+w7zzVlYj6ONFDGoNj7d/BVKxcklbBgGXhYQXsUDo+/3ixzk858m83
yWxk8OC9mc857G/7sK6oG7wUoguEEmTpiL9HFnJPGFa9v+4RVIJhP7ior5xPwMfifMxMlKqyz178
dQEvqzeO2rzGJUQoptr2yq30IA1dfF5jYEyF3i5mpJFTA7haybRmwUxIkTnyelmiHmmyhpOFUISk
dJP/Nt4n5dgJVzwLbB8T+9WZpwc3h9XLm5Ayht+hVCOWHBwsojDrLAw6o97WpN5+hL8RldvBTPFk
pR0KL0VCQ8Ghas34q2+FJBzAxX9Vpjrr5zmdJA43xSLmhcIXShjcjq2Q6L4F9ZnZoVIRCfR8H4wI
WQhtkHNjgCO1FuVmeCqYNGiTa4CpqnSFJmOOhH3v0heq0072u45+H5rJ64Ef/kXr0Q8c+c/2Kg8Q
TfPT+OUBWRTBrr9DmkSip/iN+cqjY2RQESUliunJnKiWT6q/J7KOoc9XtTMWetdEIeRWchlLWRFj
OhOEx+CbPKamVrQYKRt8Lces9BEHLF+R2yMwiE+F3kYvqTc2NpBaQDEfKyrRppklIsVIopaF+JYW
t0x3/YK91ccky61Qiui4ch60uC04B+eogzXN5gWsVsbzXQsFDAdwGq/sQ2P/QCkJSC8OsElIdgSs
4oq0qhSzBkQjUV0wXsfoAybskh1w+0eFTyfGNXbG4KNPSwzP+yhe0OnpPx6Xi0sEXIXNXZ7pLag9
OfSxZcs4vlabwWeEMng4SYtx5UyyHcqpzQ9TMa1MlVkSiI0rOdG5a/WvKAvKYGCeV3ltSUOT+0VZ
2dk7iQ5ZTTlBJXwWjhW+C+8v4BZyEdvFzjQ29mCQyxmSDJlvEdBkbGXEiTITQ2h3PNUKoqNZJYvd
kWC8vxmW1Mi4tkUhRZRcQ/zIp+DeGnKN3ENnro4M6M+l4lnIinUzXaZTolCWqn4hUNDMWzr13Fw+
phhFJpTV+LGVDIUvJz7eRt65AooOUPZienNPxvaIKOUogMOANBXm5XvAVH/3/HeaQjYVlQTf4XfW
0Wa9zZ4EWHk5P1y+B942l2N7qRcWbFoRMccmBLaa8t03xtLDP0koDGNdpOlpkm6ofdU2mxelWmJu
RYWBdC2/KQuYPU2Ncahixqeeeo0PsZBw6L9LXT9ChwQJpGHuVqXiQ0ZhjGBqEQ1BTFFfwTTaY/Hv
BEpHQ02495oLMqx1yYC66VPvIzrCvoG1te4XA6L4O39JMDXDE7f/1ilsNA92TOgOQ6p9+y8NRz2Z
77oAB3yKOD03naFAAunPInrIWMkM+wtBUe37YHVJiPVa9KJfi/qHN+rsggu72AYddEZqU4jnhRK4
n0XvydICHhofzyj2pImTTCdXQVwtoJm5xxSWGvsNxFG6krrFEJUR/j+8n58LtDEFkneJehvnlDCk
aminLTuk6hkYH3EOO+aJ00m95hodhR3ekwpvv8n1Hyp1iNDjuy8svPKhYDLn0/SZ71BlG42bMPIj
Ob1AkOUGQXLXAsb1ZpT5vZBZFutp0G7//Thz+zQEyS/bvq30kPLLtBdhsu7paAhlL/APHTs2gN5S
AcbD+LK/XhrAjVqycZqBqvVFsTSH+JvwfxtRfLRRdCrXAn1RIXGXQf5CgdqrI19c92wQNsJibAny
zmUh2D5wksDHm/e3Q/JvSGuHiUwaKnj9PUScGc3pCv3KBmSO32Am5QL6Mlyut0kiltbyYQdcQJga
+WYu4EW9K9mj1bHm/pVC/DESIKO+HJEr3QlKDyifJTI5qzH/GvOkQyhfPx02LULSJeWTIUItWKDt
Q6bvsdBW7oqHfWnkKoIyG+hKhjRKcaLiQLUVHOw7viwuPG32XhqD9UF2hXKuDspU1Jal2UCh+siI
oAmHTUx9E6V26hOsz1NcPJDAtTJ6vHJlYt//2SYb4XIdzvD6sQJy5kISvzhmb+w3ESMOEaYEIMpB
RkubdPtRSmdIvCoH78+6pcoGCScqg/qO2FoNwZ2qey5xdeD9MNq8I6wlwDLXUcIsvyw22zSW67Ht
kZDBcrh52ClsdiwNZicVrn+A/XpxYFin/u6eZJ+P9HleOzmImGFWBVNbT0R5i6CE+53LcrFS7FMl
NTuOVOj8QELnv8p5EcMa2YS+rd617UfSNjxR+Q/Fq2CYsgEKjsW1YiOa0sJ4/Y2H3i+/fmJ1MWtq
wUUKvHclHSPSGQLAyM+x0GwvMhj9RTdh9Xf9y6B25QEW6vO62ByMh54krquwFVf7EvwdKnWFDu0H
dp3v6axdfNc0ScJF048PYuUnc9H/FM4/bWVfuCbD7IpV3Pzs5/l6bLuJ/wIt7u8DQ8FIvpCoB0TY
4aQLHwR8eaHFBJUCoCwlkxdFOmowWHfrznMphg0YAQjCfMhYZx+LLHptLZSy9nN1N/o5XqIN0ZMD
16XfdQ/h96FcXqS9g9tvgmWXzF9kZX5EXzPTGXGNlI2Ox3SXRMEBxpF8CuaOGYSoREBxRmbIZh1l
hUjtnVcvzlg1292x4gmyK3Rukhe6lPPOkWMk0VngntLTdgkeFvsXzQKD+vHoH0GA/agsWJARvi1D
9L0KA9GLerxWov99ZmERQKW8Ig7su3WNxTCMH6U3K9gLooXC9uqx1NKmGXjoAuvXlqDjCx8x6hHx
czmuREkakewRai71r1CLchcH3dkhw/pGFBiLSo8jaNC4oYa3XJuWfzIxq+zWUU1FK1ROvZBCZZ57
GKpGB/2IDn5iDawVbFNWVS+nk9TPY0StGxwD/smNGl3kH0gqQMnG6oMuK372KH+jQ/EFp2xMfxkq
GDTlT55zUYfKHIumfkSqQNDrapZ8Hx5rLI0KgpKQjMusT5vQADFY4QxhNxcpo4c7oolB9q3yFBji
Sz1arIKQRrNOFf+XUCvglzEcPGlf/jp66P13XR6sQ+OhFZ31RsQcQRNXN+uGf/D/wpDK13iccFYN
UR9AtIICvehS1DvDPLz26yWgL14PRYPAO3tMFY8BSd5iPSwScAYi297k02iVRYXMDcrGAB8/atTm
LT8qq2bUJHa6Prukky32EAIKQGT+PqUuWfk7zbdbwfBHcM4EAlJW7Gt5qwsS26/3kem+GIh9dOLh
AASgaGB8b6qlW0CxjQ5Dhl4YzM2sdDYQyBxrO6hZWfTmEs9Xujf16x3dMQH9cvcN0aAGsyzRHB9F
zneiXvSGyR5RZue9vuHRbfEkDUCYPeTm8BiyWZczcjmc30IzAbq7YJO6Nmt3aUYcQKrgFSUfnzZr
ppz0m91zEM7wVYe130yFtXCZSQUpnRoZtBF0STFrXQheDvDWWkuCyslMS8TW7scKovQt3u0FR+QJ
tqh7C9fGjiWlwSD2/od2VdDhJ7akZjCpUQiH7OL9QeOKYVLN1T/RqmiAVaO0t5vHrdR4MhuyjIcw
a1nGz/En768AAKnZDdjOiOpYALpBUIzXVZFgFsEtHsj/yUfF+JNJvGNVCtdYN3ZxX5c/r2BaG1oO
9lfriJo3PMO0qThGG3YCpWEWoHfnyRaBN2lWYvCY6LHVC0d0repwpSinhZGzfRASa7Kv0x0tCZYa
LF/P523qteLhTLiVgaXugoqG9ljIGKOfm7szBmJ7wNct6tJl8Ktc21QFeU0UbHhrRpf/qmOOEgot
T+gdvCiN29JhLjjubTnGapahVxtgwDbzzcT/lz8e88tDDs9xW1M6QLuBis/xiguWDxTj9DiiPLNr
l/FiYGTl2fUC2hMhed51QTYy0dvdTG0Mlcp7A1DqpkICQQ69aNTBTlwfp5TaLukIICtsijA/sV+l
U/ZwGlkvHM5oM39fg85QERfB3J7LH9F66mqTP7OTAzW5T9HHPNFYzs6UT7S+aCHzNTSZi7lgE0ON
ie6Ds5JZV0pMENiROsSYJ6+W74iiWnUsoFAmNghGDU87yj6BkFoHL9C+XnPW902TubRSsenhNOgH
MzaREJB4ANg1LiQ2dL3inKRUBSDfGjfHl1A0qqwmhQ1xJLmuVWYNXYMA6nmnihUImV3rxHCeAkLO
ShXSycaiwilmGO2MLzKvz1uYh28pBmlTGfdFLqVcQtVOtdpYxA+mY37ijCwb1EeJRkJwKX7L26Cx
KY2KMfwvSz3CduEPi7/IK2F95tRyyPLo2223wJdUM/TW50E6/YmXbcbBTOuexa5Hz+prtG44GPeC
wFTZ3E4ovvQqLqLS0StpbsYaK9Q4wIJbu6ARofDr22QPom8PwJKPoYbeGQC4N8pdPqdXsOx5tFX/
FcDs7aDBQr40MhOh1l6gR1qtjtZJf03dDykcDS9IW8mlxApCEdCASI9+6vuNHOgUKK0rCkQcd38y
hLwrJQ/BIomWjAIDRqwM7mYsVoikkVCfLCGn0kXhmK7bSONwr8Mv0FylkJITOxtQmWR/FLKhtK5s
NZtcxB7bzbN8zL0uj6eY+xR9ghH16bwoW/oJFuECrhHkVB2i/D4iKwWaY3lDSY8di4MAVpEGJcEN
/+Ss9rLGzyIgWJDjROGgdJbJwbvVYvKN+Da5QI26RZDt7KwY7Qq0GJLR99emWZMNVJ8PIRy4bRkI
b8ahtOX9WOYN0HQbd1AQHP8WUtHKAHg4FBkMRf32ao5dW/chsAwuL5K29K4yt8rYEwD7V8XtIOAA
ZmeG+Tk+gQlA++cZlk+kr61TdVyh7geedP5dnADodj5BSK9Uj14YBtcAY3+QyJ55TrLsdeIhzWFL
K+xj+fYYlyoIWhnpUn+k+Rlx+4xUVRRUWl8SepAY9Ih814zzP8A567oLwQNaR6IWJvCkEibTVScl
3iv57DuEQvtd9tZSpr4g2wC58FcmyWk3p57gx34lhZKb5nPS/cjFyecTYQkjuSpmdO0nBy+7zUwO
wrHW5n8mRV0DQFbswIUZbsKkvNcM6cKajJCZyUr5+ZAK67hHA+S/4kE/I87fZ2vNPIbjL/ZVHohk
IdOKRu/m44vZ0DvtFfnf8llgOn1Sz6FzpQ4KQcDWqiYyutEjOZw+0aOM0UKkH9RQXCeMLZGLofpg
BuxGCRya9DyYtzolQq4NexvCnzCmwPyLTRUq6nsGmn0utcCRDgQ9ROpGgNl+q1yjk40ahryrBZrI
ZYBrnTLPVkWLTHS/DDYp/UliPeQHAcpmVoQYXzdgdrqmxMjkxYsFUwRYOEiEmMVmESUuGSDqosms
F4UEnCN+RjyQo3fGyLnuaRoMOfWyKli67+aE34sEAn35710ucXk0exCpBngU0+9QbN39bSvtf/42
95OZbGimaXXi2FXyS28CU5igfaOkRS7LGm6pfpRMND16b5lQTWFB8uf3cbjNiQeR7DxhNpImu1EV
ykYuSCI7jCVghW3/lyByGrXEeIQTSNBMQdfF2JuDVnej1HGQMi1h/26IGlEfhyxMWmETjqL7ZurW
oPl8498C9xOqGp47qAWWJ7DrhG/j8jLb8kmjdZteeskDM7UwH+F8D7IqVqF5vyCoRwwWCdVEkueZ
OuZWZMv9QgUbQv1wfPXvwG8/DwBMJvoZtX3Uh0MSgYA2ZM/LWyv9ZEisFRTfi9CZqEWLaHUTMV8k
JKMT0dfDb5K4sK0vSGUUQPX16BUITcEo0RzF9BXuGgi0guG+QBBmqX0iXT3rhiTNG0Vs8mboecwn
MZI4VF9cAbl92SNvhzKVNR50Hc2CyxXDfvVeG4os9ADtJKY5cExQ237DF9/umKdko9BTuYvBbtZo
vGA6L9h/8XDnpTYj8eBwEN3mJ8cnjz3aBDorZwlRC53vl4ia7RrCPy8MzA29zqiu/aFII26Ht6IM
qBJz1HXQS3Q4nTAPdaB7ha5rSRg/lGSb6jZjwr2CVqrIHnZcXtWlQtqM/rYUiik+8l3auDgD1lNr
t1Rx7gbnSG/QQ+Gh2NIVXFeEkwUyYBLF7zt3RlCTeZMSyMNN5NLC9w0+yL/3nSh3OSYYNJq7/foQ
yeytKJVmBrNx8v1SqQdQ5G66QURt2I+8C/t2RCd4G03pHF00TQgRtbtU7C2KWjR8jq5Dhqk/bC+C
gVhJrhRqifwpZdzy5cXzlQ1YHFnrIq3l7Q2KkgDNIWaRpCilCwdCVjjfb9qfqtirI5Z2cAWROoJh
BGeYvUztsnBJ9ZTnBPU2FJvGhfjGiTdb4SFJJeoillr3CeAx6E7CgVdLJTBe2LhABaRUSedf3rtX
Qj2rmn4L5OfKeYe+0t+9TenUyeerLfrKegpayvtT9AEVV5UHZrRDR+zTBywirMxW6nRUGhreOWp5
J+Fihizy7e3e7FQuEM3WqqT6cdagghEBtPS99+44nBSYOAY3QdJlJFl7zpj+vRGBP3VnwhWHCaK+
Vooz4Lh1wBPMpWT0Juud6Zqb3Kl2eWB4TmRabBK87NAZ+ftVS2gHR5dZWG4sOMsSjxRzcidLjGSb
/ZifrdPHJr/QcRJmIuTXJDojCJP8VwoFiU9A9Xp2YRUuz97g2Dksa7f36aXeZ9zxIUgMWlKDbOFn
S/VQufV6zvlTDEyr6TlDxdWzpYjmYNRvXUZNxdI/jRiefUAkIog3tCCPegvxfftZJDJBJXQ0gBm4
1TZj+Ua+XKyf+ZCtRN2xckNN5Y1ChLwWHk8lg7rmk3twaP1F05N43hFDL/enN5oEKFOMfhJJ7BT9
1/3CLUBtwFVZVyBfZp91RerhsY4l/8wbwxL3u6aVFEbFu7WJYoTOJEHGp45RPTEH3u0iDH2dtH3B
SOANTVEgTBOiay90bGBvpidokDPf9jDOPhVsqDh6NXCkLaZBOBcr9VM+NT8V6p6wvmP1MuWZXnaI
4cGvCMOuy0f7TU0K6jyLsTPhaVkSerC7JOwEze3zS0uPw5Ykbg2wlctPTU2qTbE2TOzJzn8MIYyp
CwhRsIscLVO/2vPgIPhoqSQADeGmqM6hki7EAXKBJD5vYkDY4Lgilsc4cczYs8BBt0li5ZpTUSVD
zA5gLFSbNW4YnTlV4pVlVUzHUwRbbAb8/bto7B/BAviJytNpzN33B3Y/LIOwWEw0aNR2KSc8ATRp
UI1i5QkDNBzJpBs+ietRcZHeEzBS0eOH4jvAr1dGhISgfAAD5UG0CZc20PtyQGsllopoiShvNlEQ
LeyPDbVDyZ6Xz1+Y0GRHrprvxu9cv5n3xCQHjHW5ewpekNwnM926R8KZdVMtOELKtaZNPPlp+6/5
WWm3psYMw/Yu0aOrOEa2fS1Pdm+xBXoIFZFn/TS1yFtQqNL7Qn/8LJzLY5NawdjRaQgsOuXweCX2
lx9G3MiHPqglljhWoXIEznCMoTQAScqPwZyCVxztiC5b9AaPDeaXFXVRd3Ee2KLtsOQLgbP0xkxS
j806Joy0Wnh5V775vKrAaYKRt3p9gdpoSD12RmTjg3C6a/DE4kGZKYwVM6RXj2VvlwPkM38vOvcE
qEQJMAjjLtTn+1QStZliazo9TXSZBs0ILYcc+/FjUTO1zo4I8cdUjf8bOhO+5xD6+edBLmI5Ydj3
KpbFruzeR6ygE6TY0n3GQ0bmGN24XJj1+6Oz1vUiMUf91FY+i+xLv//HPJUTSXMMaYOFtctUTN1u
jgTZOQgsPDir9sBiRAX4czh/nesRfqx+CrcaoPV0KThivcdYWMZWqEPNBVBAjmihDwpXidqcmZGa
uzxO04GtAGbXZXkqNxgnwo5soK6qr9YLfT3SlfnPlioX5zHIQOMit2unUscu+FhoHjf0jUxE7NM4
YHg0cVvIHPcX5J0P07NfxiCBBDGjxkIAcgXbqOuspFwibvfx5pU27r4KXmfkSrofolKC3oUjJUFH
jOQjAFC5wb8IK/zWE9Yb8c5UfZCgIqmvzZO7AP7RiXlUmZOuYUGj4uyWa5/99Li7lnmOOwJAIREA
1i5VAqE6Sj59aU0gu8PsA7jPuCjm1ebauyN+YCqJQQCn7sbv2EXr3As2/1VD44ygjnCvM8/SrifE
myfy9FFYg60U4SLvh7KOdbiAc0Li31cbcB93eZopyT1IXR9KBd+r3z5sSPNJllsqyjuohIRRUDBr
QZl9Ay7vw0OR2blQx48N45y4HMTz5iDYixT1w07iPnEORMa3Z0rmnrLFEj07M/GhuWsyY4PX26rv
FAi0nForGIuaOIFwU+Dc5DAs52bS53UD8NnLHh1CXQxAlShFFBbSxJqaMQ1onlnbrECDNeuEqBSJ
JJ1kK5ta4AlLe2J8asXcl6asKAZcDfFSLENYSE4zuLWdPROJAOt0A5ospUWHOeuFxpf3p7TBpBlq
rt1LdtfiB6Lnl6QJeIvSOp2XHLXWDlPpFjZxuxdTS2xkF3QUJ28XH03yVA2d0X2fdQ5SjCaAoKhx
heM8o3uivzBIYuDCX0mvVlsx+mJuCUsJt5YtVcVceK9EPfuNeta0ovt1gDBHoj8HVh4PB2TD9v37
JZDDh3X7jEvb4o3uCSY7HJCD2st6pRGKuR/Y6bWGofS4p8MDSe2YDzKSk/Jx/vTFsuqAamZQ0EvO
z2GFterlptZxWZS7PyCr0hxgrWUS7DfCN7rBn/i3lLHyNgy/g+77FuDl7vKpgFOnYNfPN6F3h56u
crzHXNbSxLIRv3iMLAElbm0qJmIAeIH0or+C8rnV9xxe4G+ywxwUXTdXemUBpY69bKEsrJbkwB2L
K7XZvupZz4edQ2IfLKEBYmkAGNEfq8Zacr7Wu098IuuHrGcxaLpHDS/yo+akK0GDNypCObbEi7Ag
xX8NKMDU4eVNYKLdSJ8kImIW4JFfNd2rggGgSw+xYXaw/KDHeTRZgR95EJdVMbYZ3KxqmKRwbIxu
IxRi86HFEb2RrZOb+uuMpcCXgpd04sKSShDtc70I3kHW/AJKX2XpF6T3538vOTPyKoRF6HD50Ez+
v02oxnS1ORy95A4gY4+W6FGoyTNWIDH3Vki7bYwLV7iu1ZKZ9RiHNaWdbN4jHarqfVl+4+QwMpkM
7FrHrxu5cUR8biY0hpo/cHKQ5jKiTidFPEPmS5EI5HsO/CX8fiY1x/EjMxY6yrYrHX5Aqu3+5PN8
8cqQVVqjTsZXltS0Qq8BRfci+/ntmJGRctAXcw8WGuWqCS7p1qjJG/SzwP1WYnlRtktN7jS609nI
UpjWDtkCKnWsu5pvz6sPFEA8eLz6s/kOt/wNpbd/eXpT2MH9QSkajje+xKjMQFfxDdP7bYOEoHEU
ErrVtlp/3+kECiHEWL50h/AxVt17q/ZVzzOJExXmviilYOgEnv4R+S57E5LD5Wzddn2LY8Zwhib0
iGkoBErdNyF5EF4H++zEJdHMDOgD8mu2BpOPnqTEgedGQJu5zmbOOU3kZMBCtFwBnXBzOlWmjQf3
B5rBtAZOy3dr7C39eGVFGV81nPbWG4/au1xIlvWWPg4bmJLIFF0aQ1CpVKKIBRYeBSo6ju0aQKwk
ySWElS/qyfc/OdXKPxE20XRl1Xud5zQ2ZH49/9O/AyPlsNE7QTUbpKLVkzA7On9+Tq6M8JwS88ER
cSpFX93v+b9rf538KCBRj5MuJTQHsxO0iQrCuZc4nMSvKZrtnLtab7+XjEZMwW72eHSSvq/BPHDV
p7p0F/zTvquRSLByKgUnu/dXCYTRuGa8YMzz9D8rkXO5iCOZ6Ymq9QJ61inlAlpnlf2zgi9MXlB2
zpf3mHhG+bxL9aZQTrVE/QOSAFXfsbkMRVIM7e8e1UD/HtiS6lRL0g3gO7apP4Mh3YZkymv8BpiH
JMe0ehopLrm9AqTnqSGTe3P9S7n+upW3Sy3AtfGflaWwb1WLR/mnlw/jwDtIkA7Fk85/w6sDJ4BH
WPBkP7Vz1++2H/j2FCYtNaUOanc3osnZB8VvSKsLwq38rRFFdZHgK27EfRaqRE8d+UCCTl/US+ZR
8/PaKCV80zfBTqfLIVrvU81U0uxbEPIs3JLt0xrsb16VvLQic+Pd1OD0jYz1UY0FOvhBFOVeG0le
XwkjqayeP6irXlA0frXuHUi3EYY+8wjvjF8FXA41PrLZLesLUZDolUWv+ISjDXNTv+wcS14kvExo
2o+q1Fk0Gug+qVpi1QERqVxchPne3t+o4JGoZzA44Dya/55NbYjDcItcev+zk8RxLF9P9kVoEXef
cggf6mMX99jTcT8puKcDPCBEYvBVgg7EWCj7dUhx0k2coosXsfD7QMdOV2NQNNIUm1xzmVyZ8Nhl
C9NeNaf4KjHknWKFwGMj2mkBtUAu/6kVr8TXCg6v79XX6VjrHW9YAQHODzY5IvDODstjE2hns9aB
/uOCh4MvdLm+KE4i1jS6rKQk6dS8F+esE6kW2ffQh52WkRLAqdWROKy51X8Ai45+mcvNjlBG2543
bJySQDO5UZ+PgGRdlqz8nFPv/KuTff29on87bJei4F2J6PU60Kia7ooiK0O3d03Rh2x16fqEK18A
IdXEn85/RtjDsj9O4v/gQC/Gn+PUTwNRF1zPk7k+13BhrcH2aZJveYtxDlcA/E9Det9LhEhvGIGj
YVqMDhCPmeBJnP+ZujHLR0kM6p7XfBXNuoIYPiQoKyUUSeenzg9TKxI+VEznImGcoKtsqT856FyE
CftKX2ODsu59PJZFb+5VQ0z0GtwGEiNzsShKRl6yjps4vuLDoplFCUgVZfNkh3FQvb6nECbduXvq
1/CyJaO//2jPkO/AGhDq+75xrsCe+TWTevaz6uk0jtN2uZJt0RPruAIT97G8BjXB+gk6rlYlNyGc
wsFiTtmwfTBJN/QNwWuPrnYl7pAhjp1iBkvLQR4miLsmmMFugG2qYtGkgkavgLxoDxIqhIfbkfj+
i3+foaGWYHaqXtNC+wKZUsqmygRCd2SUB+Qp89D42x+oDDIctKixmzzNFwhqVWuK8816NRBqEZ5e
aw1tK1yW0zDjWdCD10yjfDShzydITHrrlmbBpMVHIuSAGbLwODvt7klVhKNNw05c7a5D3FNQWTNd
MlpQKWuODI/bYxr6c8eI97XivLfsFROukr0jq57znxFlNiJT9YXQdg66c73AgdL8sf9MWuYEJP3W
Nkou71rjSQVOiGXnTFaBCZLOe/j50B68StRLFbnfl2AauoeqGDsmKkAhQLrLAF+BoHXvY+MJCqKI
hb+2kAhvB7Jt95ELXGyeR/lSV9g2H6Zj/cLH8qjswef+q7jMRcE57FQertv/+wmvzncloKignkhJ
QipK3egurTB79t1uTFTATgAGbOTuP8UbSjMYtSd71fXPifCgas7nqaRb4bktfb6c5VwDH1lveuff
fE8AB29dSLXkMWQNzCLnKpX2IZpvXxvyzYY10IQtmNmCoDulTIbmJ9bce7J1oPG9j59SJnVFaH9z
uZ9WFreKreRN0byBBf1rzxl4POAF0ZN9T8g+8yH0kLdd5ogGC+RszHLO7N5p2iznutCFgRhUJenY
0HAEBVcJWnyPH888lhOftaKqETcGY7boku9dWb93r07r0llL611mCMhONxTtk+Dnf4uWDy+KMPyW
0VCk27PfDl06nPpdGNTUo0ZxIhWQqVO//d17mmsHuYmsF8eTrRAyPJ2F7oGMYMuuAsG1ADOIW3Qo
uFkNjraIu6nPZM8hbWbPoeSz9gFkyLxomoqu8ZhJ25IiP/wJRDYjNnzODPia7HEx/h6e4CfvgxL+
dxoyK+aicUAK3n4jzvbC44F4i+p5ekZ+O8CA3ku0cXBasNGRaUB4f1varLB5A0DbXUhtAhzjmZ7v
sw9WZYqQ5vY/Bzrf3rACNkydc8I876xJzsiwx+oOavXwDc2fPHNj7nq4S4nlpnjsWooL3gT4zm68
Oj8ZHn+Bzq1jrpVFro4ExyJhQwyD6fxuw5HEFSWMsyeli+hL4bvLme2ypfbqshYPd15Sri7Yq/6X
6bVdzpw2sTBfzdrj/0F8I+9oWN8ombxk2mIZs2iN+goPG9XpETRNRLoR8F71ztTXJg8t7LO/BeAP
UYkLCU9slnXM2UYMoYskr0Z8P1Y58RLJwwbPI/3Ow85eFQPUldCIW6tJEQXhfzvsCxhJQLCc1Zpg
OmyprDlJ6OGre/WnuXNkjjWTssfgJqnN9i3y4q6TcV2AlRDQ6jqY1y34tuyd/XhnI+RnQNFwcDa+
9NzAyK9wQiEEfEPkBmk2Mj0F8/6ksvijY6OOyWSktJFeEMa6CPN4l1oGiw4+8dsg+NtQdkkOwUaD
G5w6aWpVfLoWNZ651jCY6wxAHgIynaLWqX8kozY+1tcdb5AqTMLJaWUiLc0MA16mfzsUvUDdZBMy
OpeTSQBo5Ke7jdKEZG4HK90TZft7N0+KPqkHeZW/CGAUane0u2xFYzi5jZ9UFrD4z7xCDw1GDo/J
6CFCmpDlo9g05awrk/fC/dQHhaiCVQIAwIfmXFajM7p2qbdJj201H+uYiIZ10GpadNCjiVTcRzBY
KEq9yoZ+sk5ksuww4QkIY/yEz/zHJcd0DKjyqui9h4lmKsefLMJne2sk51EIVPZ2Vb00aNj82T9P
n7qEETpWHGaUVr5dBu3t7aL2kXT7beoKyaUYoZ7NNRXuh72pQV7RsZRLb9ox0Ba2qdq3xkWoqElS
RXDGfRh5IeTlsjhaAKfzwGpCx13pOp+T30OeizctmWXioFzEmxohyxsaBX6wqO4xkkD+hXgRB3J8
wQFsb6b/ox4oB2Eq3AqLcOLYtvwpiqADW2MDFQfKyECYQFoFJuOk4LPveHbLQYVUOsDevVg+OQ47
fUSxEkI+W2Iqzhu5t7M7Z9pS88rYd6zCrjbVmDziAR++y/4YsAAgVr5q8qivaFAYsEsNlT8se6pb
L4lIHV/bUdmo9zKUNW8iJi13lB4hBLBiWXHChqYacHG+NJhrbK4lqRe98f4+x6Uo7EQOtNlXBv0N
UiAt5RQJddvnPO/CdQhgjf/nie8srGus/i1uteBtD0Mpyg/PQc/sBUUTs6E1ZVdWdgEn4CcJMU2O
iLlM/ChHqNCMoBjnJkj2y3ZCGA7M589Qp49GRIQ2QesA6/a2afRMpWVn9MUwyolJ41q21UrXl2Ib
DITlMuEzi0LvYzxBFLzFMUWzo7jgqDk3NQKcMYpIXhoTuxiX7yYF/oSJARVaSP8Oz4+RwhNBZ6ki
nw9Ahp8FYCmi7SyE9WOEmoBq65QobI6EOldHiSfgDqBLHsEUqOa2iGa4fgpXjqFYAD28AeQevDUx
EKdujOBkIEY1omsDpAsw4WrBFRL7eEbhpMyLnYYfqsCMmH3xz0a1rOkGU+/WP5Oq99AOyJN0XVUh
3zJVyF7COshUQKClzVRiLXSNmAn++WY35zASAkx3JlvRUcW4otfzS/G+68uVhtDjAOFWYMdHdELq
sD4VsFcDahZK/p9UMEfVLUBmz1+Wr0rwDPvkWxbJ7OJqbf57n/SvX9sks+NcKV8GM2mplIKpy5bq
kGWP8eURwscnIrvO2S5KdPHVq5rUM2MoqlRj7CCrGiD+emSC/VgVyWmS9cxKU44Gh/1KR0kzVIye
RSr4vgdSe4BF39Iv90FKs3hLAJ0KxMBjUcWLDHHp7sLVdTOUU8+tZT94ivcixkTMbYGkZnuf24UZ
mq/J5AYj+ZPlLkViOSgyKeDd3VIrP/LoBXYMAwcciCEAobH1LQWBwyFOYe6xKlD1bUlOUlvZlF3G
cvfhxdCK1oOmWNfqziIE4de7Sfzoxi/uKJPXh/c+q4q2li/gx89x3BsbSAByMhCIuCWCrf3gFg+L
j8UjL/XHj2DAFCfQ32LxG7ulYuw0Si7Yvq3+P0RFwRkFqhFLn6xRUIA9pMjF8VO5MMVQrtrDpg4p
qDVH3gCPva6dynT8ZLnDSi/vLRRI/VQdjb7qqR60WAhQnyU82Gd62KwKRw0VFzorgJzzs4/HJO6V
uhMt65b5JGbO7RVgSNN1dcDXyTQlJ/w1ReG6xsN/H7N0styNQ8bKWk0gEdE1f7vvvCvVv+JvUutw
Ker/XlRjX6k0tOH2lp9X+r7/M5Wv8GXc/cFORhyf4jfeoWlE6OvBMUhTZL52kc1ZLCbAErk/QSkl
FfD2U3KFUEbGKsceoOv949gSJdfZRL4aACo7Yp8OXv5hyY16A3LY4kDuRIPO5YSx+RGDzaj18pVk
70xhzQIykmxHsYsKXn+pDCqyfzGpHUl5KWclB9GfhZoC721Z0OPlgMsFuh40UjCnk3HFAgRlFACH
2fYtNxJLEiWDQ4S8ZW6EJxE0czE/2VhrPIRaBCFFYhLGoV1Qo6Xe9/wZYPNSj+3P26gtOLQ+/qpS
0mEgcVQBB5uBdpMkUvsVakAFLUGWPf2aifuQIabYv/iMT0nGgQGDj2hVrXIfPtT5P9I/y/v0i6g8
QyewOJ+HvQS5ACGqIVhuyefQh5YDsNtgSg5Z5i63OfjoaayMVVXWt3qkVKEnsy5GRqs4HNAnq947
fyZ4GZu0u5dkXSGKQrBlFKwHKDKY38hEIXIm2OP7GOg0wMJrEosopRds9OE2l9mdl3CTQlK4kjYb
iO0JsYsDJ+wIarLGp0m/onhXctOUEk4tIExVoexkPfdOoVoonKwVrtpP06NAquGlcLOaq7jpbzHe
3NFhE9ndoQz3DImQPmCo1h4lM+FKXky4/xinO2wNqYqfFWrgCutiwpC1RGwMeqszWPBzfv3s3rFn
e/QdSY0YamYLTIsEMwE9O+GQyjK3rx2R8dJpdAQn5Ar5WES93Q/GQfiGPTejzipI36hoJqPwUc5m
5rhUqd1Iapxc+fg446/Vdn7eoLR26FcQ2IXwXMKBS7GhZbHvpmdpVNYIs1H2pfr64c4xGfM8Dq/y
H8Wm16Amta3qtY3HoeP7cgW+vvWZGzbpMCHtv7hy/4yNEekBN0N8N2KxHoHLo+CpxOVrQKAKYBcc
vXI/2mG4TDXjgbcAGfmeNVHS+Gy3jJFLWFZRUKA+ltopVqaUmd/rsiW3iycyEMZMyvnjIvS9smwN
f/fBcWyyIOGKZx9arrN39Lq9ifPFs7sj7Uujn9MrFLlRaS47A6nW/K1DBWMZLpyHcbKZB8xyKHrQ
QvB9dPALPBNbautrfVjcscR2tkyQjEjJei4fH0ukZ8p9i7Ky5Ml7DHqz5OjcfVEjSOcmvINcJ9B/
s0nO6o2JK210NclU2eJ1fski3WuayRTqu3kHRRcnNsLTdAsiSaYThLqWnB8ttV7ZtlaNvsoqIudF
sVCNlLLU9gxtnt7DFup/L9ENRjVfs0TzCILrzJke/GyUmVdrYgISF99qtv0jkGRw3ggdnQ/rgKMv
/VLeMAekKl6MBqQHS3lZ1g3JV9GhvCGYQrIN/BUvQYmxBhrOMvWVo5hwwVAgAqrbDCiC3DTUp9kE
1ei3svNIu2PkRu7wszHfvp4VolYxHARZ9G/evjNaq9Ch56KWVtOP1zDUlo2kiIoTvjGDf5f2zy4q
fhe3YRmaw3Mv1TT49yVQVLH5i2pfrWcQbSBq725093luTFlSvQXZ5GmmmJDFRJprOXb/N1h864gO
UdvMds4oFtG+fqXIpNsKr3lrRlheg3gWm7WBDtwqrk/pWbAUjCH9tviDwy3SjN6CxLxNjfaVvWze
ZBvnZrUz9ro72lERjUZH+U0ggmsj6Iqwx0zH6Cc+ZMaqK7B/X+87yNI++KOfjiQ2CaCkD/WJjp73
kjsd2L9K1Gt+L/R1pDrS7A25f33ZohpoMulWjPjZhT/wAsBA1KAMgo3zczZnyAltnDVQuZdOxozl
yWPjYlG78rXe4WGIprEFZwEN9Y4TeGcyG5Tcq9YCYF3v8Y3xAk5ee71DZQTKwOQeXvMvRqsejdZu
OxN22PjIzq2rvlQCqxrk7YVQuxkxJ+ezgtW4gkMiDJ/utr3EahD79ElrbDe7Js6Pc2x3YZC3N/SZ
hkXt/QsAvp7ZWXNeYNatNZ5A/lb8WxsD324gx3BD9E7uLsIA1vizUZZBl1EFt7uQUAbta8n5eiDh
Uwgl3vnDTLfyg81uploWskBchApluilH4THU+Hx2XykFcDsTTnYkx3aC6P3mYcxwfuIc1aoX4Bgh
WfDiUTMCOsXK0C91ug41w7DI4l6LWXuRXyc/ZDEOtIsJDXWRQEvlBVuFsoQqS0F1fyvAx5yVgWdE
TFtLd9xY7haAKWpzlnlD5beW+ocBIl5rhsFGzpo3pQ73ye7ZMEC3rLAwy6DnCz5aDaisco8vyWW1
NXKNhUvA4CbERLAblAYo6Rc/z6N5JfvnDiQqF40Bou4KxHn0bxysDyZ7MmKrfVEDdU8V8LCZzKD9
yytM1FYD/bSedrgI9o/X0sgyk1BrafrDz0ZzXhy6DJsL29I9EHsIwTJ9oVimmxAXy1zLN7oXOVZ2
VmdPC6OzShmpn5rcsFzmOiNuj5nfazloG3CXR6LZBPSKLwHI+apsC/Tk81YSW1wYm0spAq20Jix6
8lgDJmb7bOO3/O+YcN1ncYVlNp8kCeq52z9ehRNPb41t++QLOFlWvOyH1ztpYfqBsHgUyjohl8bK
0oBtDE4QunPnq7kY/tMsrAMqsLpF3/8gYKIaAzX8IJ8xU+D7EMtoKB49Ke4nAL1dVz9QOsAoqeKm
UPGtWQzQw4W5uo75rTxJfOXv66F+XUSgeb4VGmc9J9Vp9G4VUngT54bcFS6OTHMy4GoXdtFjrZ1s
IDBCWecyTOEiVwmiAhXk9W4QUHUpz6I+nTsEAVDBOGDkZ0BipK3cP/yHoq5f9wTTomZbR8vytC5y
S3Q2FEQBHYkDi61uDO0KSh/1LWi71oKrSTfzofRoGHG7sE62MnxsRUyh7MvfA8im5QwBo+aMW+R9
Q9RfgbMC+gKy5W7p3xxsRgF8isi7EqmPXKACxqKL/CPs/bUEzlqW/0afkOq3MpeUaPyNY2a+rUqa
E/z2yqmGLDXlb50CdFl3i1ToM3j9q1O6hxk+dOr2UKYhJupqvYD+SuL8F84AmAHzIMzbg+V/pSpQ
14PJZH3e17yZ9X7z490ytTx37a9+s/Ss+IF52E2R4Tj7GoaRFN/IPkUEhT8RWSoOz6R2Tbtu5mBi
Eyma+LJhjh9PMnYNeKDTSB9Bc5L9a+64+VGS5FmnOOCz9ppxP6IMiJz9N+L5V3Otr07ALXOZrx3Z
6YoRVg8xJeZcBNStJHlLvHkvO1QJ/azOCp5biRylWAYGcxrc6Yvdt6gFhGVbspOuwO8sv2LNKWDn
EvPRPaTV0KHpE6ps+D8pbaNwW57Ii9PS7N1IZwtr1nEkHwReoE8PUsS0OHQhyf0fqS8GetrMm6Pb
5U6k7xCuPrPZnIphZdyoueqxLkYjZnv0hYHbGcgg+RDQQm1pNGV5S5lvC3hBqqcebRYLbtCuxm0p
TAdRjKE3h1j4bpgPDDt24WeN23DukG9wCbFKO2Osi8qdCEhQdvVZ4wicYZLiDXVdvY3uMmbPA/1T
RS3kTnJDvUXLyO+1fghdfnayf1lAg4/frqiPd64QmXuColRrHSF/7zzpBSwmh5cYcGsAXRIWTLyd
wBWqBP/668OFNKxqXgc/xDaL390xX+wCziO9ZRiwq7LlFygeDVmpiqiBPF+oinVcH9obLksVCdqc
/5BxdrjRkUGBMHHsyZkGJfa34odhHD4HWKpsuSe8xcOcHTHYeVuUunKSbMJWT9XPZY0mXXCp7HOU
0LNQN4j/nK6fE9NKmvMqgI2yAPiMQXnORbJKvJXJwb9GhyLDCz4ip/AJOZaxFSTDzKiM5TzdIJ2t
FL2xCGVrHRftKIyDUndSiGqDoDqpZPwgvPECok+288gktXuJ78VzZb+KQj5rNbfGPnfRASTMM7Y+
xC2QUhjqZtIY/ZBRvhHfPBJOxq3aakna7Qx/XR/prJPMShoXCg/1FREnpXKqeq5NcYjM+Ybe7dBw
ieoOUDedaX+HDhUxiTyDt+yi8T01kxUbgHmyvPu36wPtrqve6ht28SDkMQxKQhqYhdI+26Y3Vnda
c2O4czye6Q4l3vXFw3VnSVnn8/FmjKZJ0aDGgBbCBdQ/a9PjaQ7q6TJHE+L00ao8IuqoinuW0Ql7
4Wn9qXqdfdhEBRAPp1QYK5EbrLN/LXDLwqMklr92cUBSvzSTxv1/bLh5Ctlj2Twv2Crp9esMIVup
tpgH285EkMz4VNwtwWhog99e+uAUXWXEZpttcWdvEoN7EsjwDYa2txeDLWkG8vBpxA41dn1rIQns
QXndyvKDomb2RHgtBnMfj4e5sanjG+r5UtioIQLmjAUG0xnkHUVm6FXvnczaAQIDBm3aBS2ZivA5
Dg73y3bVjDMVVB0VwaSnYy1osUVGXw1gJeA4qblKUg/gsm3+JuBQuur1xOqH4dLb+GJ+6ma9Jman
ds/SyhnKdz6Ci8LoLN8dUzRyeUa2OQzvEJMNLSwTX3dJ3sRsEKVZ4V1GAagwc18tDmi8FkT7E2h2
UVgTf4rLJ9OAL1U/OTXEtKgy43rkyN03/1BEPFIo57KG2hgHVTuX3bUAiikkZy/Cd56Sg7XTFx7K
yDQetUblbkg62qwgIegIUWTaxjCSq2DH+npg8jPTmewZhQYs2jzW9hJ4fU7fqO6aDIEbA+o1Bzpu
1EqhemzABHIeTbY7894Phl3miZDSgswymJnNVn6Lq1vgL2kVxBlwp6NtMJBhjqO0k8UpiUK0foaV
OwXBp4t3j41ONe2fLV/BEvdA0o/o3I+ja3iq9Yzswb+o6hC7T8oAQmUSiVUhOPwcTa1Q4rcrOLvt
JipMKhMpAmDZdC6UIvyBV8yrurMMLlkM9NuS2Z7zzRCVje3BqqgiKCQE++e6d/k4/JZ56/aGw//G
RYkJQtI2IbOfWTHaKaqRhQbA/H+ik+fTg9eIkdF4SxERgHQofrRYtBaC9znDBxgTl+B1oVUdsE30
LP0LMyR2JubrUPeb91Lvin/bIEVmEiKQ2eTxroF1FxIH5u6yOEITFLxnp6XeAQ+KJSwCFnJNVVYD
ny6HQwq7xdRbWl1NH5OGt5g3p3Nhw+x3nm4BLcQ22T2aS6+hrsfwFgyPDXqVWHhp3a+QJ5LosDEZ
zLiQIL3F4q23f6azmRhu8yxhbQ5lbqV83u+pSs1XflVcyn/qs0o0sfpPBOvpQCNI6bFAk8tmVTo5
+EJCkxgn9QlhghiGeK6YkYAAG5kqOijUitk3asMWH7849g09/Q+9nhfdaQeSUPsby6sq0tIWOZNR
dQzGG3jup8BdhtM0MzAk6cuRg1QXqRKHLrqaXRMEkXzVT5onNpixWHbzqTNdl890RSC3fJW6w83U
XLqNvmETjYXSKdzRuUeM+IUguB+u2IpbnrxdRSrjixY3HNFqoJvIFvUyzJBKyHJj6FrGtAHiRtJn
s67eygEhyJ2M3SpgUitztPDQuhvm3BHLP5c/QhDhYdcLqKRuOgxQ8UD/t7NbMDVJJw5fwDJ4zHRx
5KpLxi9Qaxaz2W+IlWj+HHYGuifFheoZC4MSLllNHMim4qON9QxDMHfpWQtonsb+JFvkljd9PO0h
QX5C7Uk8my2vMGnFLHEPmT4NKS7s3K5+yHvOtMKJaMW3io05w3dKDnr9eSHRWoWBN0zUMJPJVPCK
Db2V/evG0c8NEkRa7lF4XGVl7eSFBPqvcROYTemW3DgG/V02ip55cn6pMWh+KQjlhN8sydxBKW4e
bUdspe6BWtvNY9KWLcXhRzUAFwQ8FD7wlrQyL9AD9ALuUeKnWZJN3AXk0PHqUeBRKwqgC+qOmTS1
aWG8iqHr1xWH7gzm42f6erW1lsoqPiIKPNRx1KHkmOmNA1OkH1pIdd6bDwli0SmYUNq+3Z2rLJoo
CjZ3igAiGKl2atov+O76FBDNue1zSbuKzNfj0XawKIMxNM9Aza9ih/UUOFWzuWjZCKiTqlyOGt7z
WpQ9H1Pn7T4FODZowoK5XxlZa8UkrjqKL1z4B0+MVz/1OGwEnL16NJ4r6ngGW78TNOSam6LoIIQ9
MjSRPwyfkeoin1Mw90SNpKekdymp/Ynd8WpgkNAuK0vcoW6Pj/A0KreQEJdo/8H1i8ocCUNPTryT
Qv4YY3kigtTdiMCQshMv/dm4I9G6phNjqUEiTFcQIYU5Rhg/4Vc/kjQj04iE39YiPicjuwdt3hN6
dvuwlyiriOZfy3PnnS6v7J2tphiF/fuLpaBSvJb+phAYelxH7bnYA4rNIDqHc/nQ5d7fhmZE3trw
Lh6tNJ3J35zut/oFWWZnjwB2sGbaUOFAOja8w/uef/rDPQPpwp4p69avOoYX+dlDjHPMBaPrwSdS
0qrBLrhvNDL7FRYt8BeJy/5+RvwRgYSvJzDkeV9yobA1+axp//RNyyEGls1UT6UZbDtnSYFS1Qmd
lt4l9KkghnjjsApx7ruE7clKnSftKRrGmDw75lgjjUKQ5dVobUSx6YEnFfQ1Zs2NeUzKt8etr0VJ
/H5UTQA1x4FEkgr/3BwCRSRjDUENmLfPlEITQHXRXH6Cl6rAH+ygTt1WeSqEKkq/VWoh75lPBh1a
h1ca/v8h6Tlmg4cAyUR/viSJw5tM1o5uTIPbOUmmiM+KSgCUCsEJJ3b8A/2iVn9zV96NdTOT37io
HhUVDciMI0DgIzyJb4I11eqacB7QNGH/oJy4XDh7IqaNXnFfSg8hlKBhL+T7a3RUqE/ZEuEovAaa
cqBTU89ooFQmH8Ll74hiwH7miodN1jnV2k+t1t4aA3AFcqiks898inFWcgb/KZ7hobKigFEC3c7h
XYrkp/Yczqb6bBm4dnTvKxz0XwiEFHNOm8d8QTg1K+uem4Gaw50ILeiGemAeSnJ4uf1AuYzCI0cU
7GFQN8djJ0nru2UiZkpvwPgpXIBYQ71kRgLlUic5Ug0o2m6k5fh6JKuLFPe1GTV+h7jr88O4mwuR
AYq8hVLz1876k71L0sGf24/PTZulR/2NWUdtgbL3sTpjwtedNF9WhxhcWJ5nsXVVNazd5KD1162l
eCmzbU7psC+eg7Vv8OoYfXa3ly5X+ZzSG+ch5+brprGynF0kMNhXGUXWxbGumb5bYgrmEKWVA447
IPEy3tDooR8GBL0uou0V4IDEncTw4FbI9nh5T80ipYjIMnDauvHjm4vs6S3C7DUMe6GizBfJE8DX
Dg9Im6vJKr4iM+2EFnX1hgZOsWJ1VjJmwiuSZGCKDemnqT2rcAET0Un/IepgFKJB01CdPdmhDlXx
2NoOQpd3XeHotVRoEvLoXXFxUd1tiRMXb+cw1vIuUBmutRWb2AYjTs/8ZP9ao9/7M9F1SLlGJdDK
lHiQTmiMtwQ9AoKHnEWwbyE4kjFZx5r6zJETjKcgXilKLPSau53OzvkF3pepGUnBkOyK4MiNbU9U
yFAUzAU7Pyk+HRBkX43bjKUGAtLWYc0a5+aHRlcyBEzb2SY0/XGD6XAzkmS+pJx/CPO+0jqYeYkb
XlzUfCC5lKKKzuNzt1dDBiy/Cg2cTJ3Mqvbfq3/jAxoq+0aFAfYe6WaWNleYdjEqFbYhHFm+6ReG
zhEQE/4xCaaKe8vrLursrk9AAbeE7RjbGgyFqAZJ2HYI9n83xFnJQpg0i8dj1P7CiC6Z4f5554gN
y9Hc1dHnWiDJ9SoiQyzsB/Z+onhwC5HymiOnKccfnJ0Z9tSSgWatwWWwafNt355Vpr4KxbJq33SV
Ygu0AVh+BP7wBM3MWksWxCjGcYUq0DkTcMs1ztw142ftjKBo5agpO3jKx/ap4QYtTofI/NUA80Cb
xHZyXNj46bA/Rhx5CO9IUgcRegFXurJTStQqAyF79vQZuM/F4V9vFmEKywjE+tB3Nqo/zh3EgwuE
JeBNOHPs+qdfC5mr2NPOnAwuYuU/DzPviSLwKtFl4jDTDqw2vX7yB9qe/IRSZ576WY6C7/ZgW2l6
kKRHDkrsi8d3Rg4l2ULgNDV6Y1DjbJtua45qBGhWlHHsa7emmWhK/CVPjhHbtIyW6b0HHYIJzvki
egDz5xd00A2yhztDwzeP2bHxbcgynyiDtFl8MRHNwvFABdxeo76h+lVNHnTESl/lkrN7jyXyA+rV
lowo6aHvftO+vrcxeulV/SW/tM0Y1CDkION/0adE3bPqE1GBkWzq7ZPfejIrlalhIerl2bWtrPuo
GGuh291sNikhrT60xF3f5Hf/NxCvtNcAbhSmu2yIwjQ8i2ZpUR4m2Es2qOOqNLWI8KVyOkaa87QT
AXT2gEgnB86jiBkiRqYV2WIgyX33xfwKanrVvo3RP+e+KUHWq0E37MVnGdQkWt1s5uFcUpfyA9CU
sgC7fOfl7AQJ37VGAhnewPUCTCO6j/SwC2mv8c7os0rzPYsGKkAm/FGANeZwEy2yIsBHuVNKGec+
FpM7v3bJ7GGT/xmbicrRhHGfmq+0fZ+6tJ9YxHTEgbJLo+qe/Yi2oioTz4AVIiVH778wkT83d98i
gQiJBiBMbOiz/zd7CEbQ4DF2um+Hp+Tp/LtcJljCR5B9AQXFQnIof5H6XAi2ERvi3+KfNMLu//fU
0vztFLz7HRkC+kvgkv7xQfa8ZMOhKZ8Qm6S/1dswT4xu6VabVrjw/T4pzuPGSnamDD4Ug/n7487N
AMQEM55Zi0Jzmu10FQuhIUIeP5ze2Pth+yTkIgWk0TFc+6unT1SctfkyDTQ76/jFo50F5quPTG3n
c5MoiTXmCP9qVtpNZtJCCN8nQ6eXJdcWZfw1XE0MBQUySvoLZqZ3HsjbGUazc8OssimsuZ8lkNJk
n1W/agKx5dL8G+N41EEiGk+YHIH2UlrtlBu+gIgYYJAEkiQ6Y6Y1PM7ZqRExLK5v8owJqnoFcLzZ
NIAf6iteZQ3kUE3zmpG/mXztDxYNjvf5TVQheSEKSrdPQ4KPqtIYYtftiO/HyJBJDHlRmq84+OtB
k7a99GPFLvfzpvP8hAPtnznBNbGMfP+d/BpOlUjVWmRbbUWLML6hE52jvVOdwRmnA7Pfhlf46x84
XLSdNXfO2ThLKNYs7ZdwmrJN9J/lATqPcpD706l4bBLmihm4lE9/t5kiC3mC8XsuukPRmMkTEoFL
aVSmM1QcDHzYKFFVYZeUnHu5bLcNPaQ7TB+DeWzjBnr2918YJTDtvYhmAuF2QxpUJmonm0slxClO
Wt6flI7T74YdDX35e43Hf5FVXeyRDsj9LLP7Fu4fF/UU1D6JdoGMhLw7DjOi29JCjOZgRcO05mEk
AAQArtZJO+WJW4E9FaVhYQ9DLxUh65xj/Ih1m45JREK2iHIIp5lzvy2e2eAkTppaOXz9UTERn0HG
NkwcCp8/+a7XIfomk1ceph0+D3iQN8aGSUyHVvrl7LGMDasPtcDwNw8S+XYgUOsU0+B9fXdnnhgc
KWXDt9RHR284l9PSarKYGa/nrm0MAEXqH+nWOY5+OPdfIj67T4V1GtlOtVDiIOFEe/BCwviDOd7u
G1YQjdMUZ80pZ1qhSSTjDvwPTCnLM+i0svXnkhLc3ojkES+/faWriuK1A6NDYA8adA0iRiOVMsIg
jmOmsDLOYJ1shoFwXRrvJoDX0ifV6kKMu4UagXTQFPRrO6Ttet24RbWyYOqlPZO/eMHoqywLCgdG
NFHa6CVyjmiwn1tRruWtXYpao0s5px6fJzVsbteBlHFE9X6L7hRMM09oUm8xu5IXU9gimPSyhPY9
lQSbOMzrbX/vfxVeBz40fICe1mez4rm86haAobzBSctdX9u0oQGvJdbpoWwQkVMYE39oJ7nrHYuP
j0Wo1ozOdG2gTjC0aQUcUfb/EQFUrJn3xlkvEl9LG+QvpXuOnrDAF9MeHiXq3HUbhf7330Pbuqgy
e8tdf+aF5425q2x4U873809VbCDmW0bVX3fOIYFTBR8/CLibbP9kefLjk+UswLM2nvJ3Om9r3K8/
6THm6YRpqdrzqvfSmLcAOe6lJ8zT7yWmpSjysIf8TS9G3GmwLUIaetxw4em+9Q3UF5C6mXPsMFjw
evbr9s7MP1wR1q2gdD5HImK7ePgwLwK1ugxX9ZaFCRQSv22rMFSOfDhimsAWadFXVUftd4JEhrwy
FZJvLcwzCC5CiVE405feh2fZD9VyyoaM5+xgVxlqGdfLe71EisZJHMH2hAXWTNlRq+nPVPo/E+M/
TTCulD4bUQIupbbaC3WYA3ZklfLdihjcDLHvFBDGb0JPklmjO2XnbnzahOPPDM9xwWR54Vioml9o
8Iq9tkNY+SQH23owv0qgFaMv8hO5PFrlJKBYOl8LjsiGPT03nc2llDd9ki2tuq1NXHRbG/xqIJj2
/wjjU/3fmzM+SN1xAKOWREURoyug4DiLW10md5skmoVaZ+cZ+5u3N9roJ7ftQATNjLrFTPD6nsVg
aYuU106cfxaZs0zKAHss360rA/AB9zF357LFQIjJYYay9iPbiHoWDSAYB9vPOsMX/oojes6Mpz3r
JkyUqOF5kMjnQdAs41EZD/M3ALLNgFOP5Um7dq5GaoSpqAeSWmNALjc6ji+BDh6/UFilzCuexSTr
33wO6teqXS7D2zg/iytNpSraMB3gGSN2ChwgNkawsUJCzkfKW2sdnS0jvZK6N4bepYDFIBVzP4sP
Ie0yLsDDaWSwS1Hme9hV+Sp3w0On4ULoci7A/huIAJ0oGzUjlpDZXmdd+6G0W4yCcxV2tqZfmFuG
iXQTrPaXHb9GZIcVu9iWKXAzdi8R7xFtZRXeEVK1LtGPUnNcb+KwPd3d0UFxSzsaylEtwPTX46Un
8O1as2DrY5Rhw71io5Xx0joNSQ5+M3KK5kfJYFQx0OXzGEUKq5uF3ZvlH0rc1qYlJrhKtz0Wc8zk
1c8xZzY3aJbmO1KQMxdHFfxod/PVgZ1iAeqtY/gHeYzEPhJ9gbX1yRP/yBu5XCIzgcdAm5avUbfE
742WjhwAQXVe1+t4Hv65rjWJNMWuilfeEW2TuKGA6ImEhWrbMci963NTRcpY7WHzZKi9DvwH/bjq
w4H6ct1G16JK81tnPIwh7rKX0Qj6mXkxlfzVFbbD1EGuNE1dKW4VC+t7Qao4+LXVqnbMPQkDvvEl
+DYk+Cj0p606kaMRYixAdoY/7BPgmC8V+HfpJTXD6o5o2kRu7cyHko3DtJ2+OKdPaXvbPZR5PUAd
+LxHybmg0miReZ4Hu+7z6ZL7hJfyUwat2Kxl9r1K0GCOC8BkqQGEKmGDXHUpC7ioNA7KhfqoUe1l
jnxz+LpRYJVIhXMUHD8SDZoCalOaYEfgVqU2zff/9MMqfNvhuPmdJKj3BO8pg70DJ3xaK3CFRnJs
guZPym3GAUKIbee32Kg1w1R8hIbARJGlAkM3zi1FY4eKoVOJvX3e/z0404oOXjC1KD6UhupaO23H
hepyhE7dI0VQk9DtvqbaoJp4Zsl87CTznowpQmSq8ZEN5A9GYmnaFMk7HaIkIgJTbHCf65f39mqa
6TBiWEd7B9H3W2vMWlQBGNjUqFWE5fOrTnv/NmFAivmeeDG4Qf2QupNSgn+AHmQppNwtdudtpw4/
3P4MwdOasZwliWZE/HcscCA7XqVVRb0vxvUfZtYw6+m8lqZXdI+6YknCNs3v+6tbc+OMpD2oefH4
DJhmOv2G7vUliFBHAA+q2wWLfFKOFmCMxkCohc2vzINsG82gcpdbaW8v8EQMZvDblcG4q1ukKzEq
1QgVE50tRb/jQb7p0LbqRqHkWQ/gUo9XydE4kTDpFhKwL/DnJq1u8h11+IQyvDYjtT3VdSXZa7+d
WZW34c5lGL0m7MFgCe619mfLaG+WvbmtvmzgUAlrtdDzNnXPp5kFPqFFWzlx8gO5NTiDn6mp+Xdt
D2oulFi52fgsvBkiFIsYCVNL1MDB02nBR5o8DJwP2/KkDtgBZFUAwadwfM5hYMbECWJzhTcil2ZV
1CjpptOsCt7VHhJaM5OU9tcx8C7+ahotkg/Fmm2Ul0jfES8Qk36enngvxQ4ORtBQKfKcdGWVE+UB
nHQfvaGnbaD/l/8/muWNb0E74ugfmHs2FlvvErOHya5D0injECn0wFrKiq2MWmhUtoc3+TLSQU+5
X/7wiSoaVVTUnjw4A8we7jY0fLKDrHOh7tzXXLVq9vla2szz5nnGLSwx2k+HG+yu45/rUgCwlQN/
puoCfINDHRowOphnIYrGWGzM2AJLAFYlUR+aH0Fje2wj4oCyvVeAXmWFqYx79/Jq2Z633u70q61n
cJ6Og+K0Gn3K3UzA9a6RYN5lo4lgVF9UAAZtRBWe0lX+Hyxr4LpopEgqZS0Z798toloMceLXC28j
HO5t/qUFdSk+bvJDdjF4MSx5yRcMTiQRmnJIehyzkZBWbSJbtqdE9sS6qOxC+lL3nJH+E0xCZ8iP
p0xlNfVOYi6BIhVW99v5vb2wWip5JnIUVbZ/DU7ypsxR3OwJ5P4V1uoUx2bE/khjfgAcPf3z0ZYu
0rHRzf+2efV07509T5rdXr2YwmziSmjAHaZ+2yidMF1AWY90b/BZVqxm/E+XHnFkdihrsC0nkVVG
k00rk/zsVmk3+/HXdEaJCtH19gEVjiCwZtFMldjTJfciGrI9qfudRwmmd1MbQ1XmPz3BTIHDCmzM
p8JEmD2gfoUWPgiHgPV6I+xKnEAr/MY5Q2AGWDhQzQbqViLhxRl0tkpx//Xw8fLYPTZavUa3NOxf
IFtcbSBJNMtctC5L0ZYzsk71MaSYuYqvK5phUPVYI7c9hKScu3M5KAUTkUhNXKfmkYz3gryZYzGL
ZWV/aLpGLEDF5cEabZrU2XLUdp6mdAzRJt00ijNdAuLxepK2lYkdYiheIT4iBjcAEWn+z/rOQWY4
YCBJ36SfrZwprtzSZQWiXzMWZv1wWzfDVJCRFfmJBZFz7qj4s1Ob1sLDrT8kEBNhv7Db6nFmMLTO
/kQUO75UxxR7uV44uPc4yCFXGt4ZENKK+eF7K7cdypBohuRnU0wH2cZf/OF8XUvnLDDm1oI1GYTn
eiUMagO2pKq1GngqjVqRXFl3/hIBSko8uzsqffVCKYIbsMLemyfC0Q2d++Rl991Ol5QLKKzRLXti
oam6x8rCQjZbr+0cXjwjhU5I6d/5ZtC35+1edLRITold4ikwDS0xMdhoKswOGn6RojWnHwq/hb5C
DAKeu83GDl1DZaHy9AuIbUhjC5HOKR+4DzPlR2j9GwmpyDZYW2N6tFI5GelIJbTvrDTxvh8ZEHq7
1iH9fdKClgQcjz95jOwQRfvcLQLKzAkk9Eus4oRhzYh7bxJ4e045JhOCTHvPio+d+PG7v1EYeeau
AAc5nCHdFKG3ZxxVStMd4wwsSxnDmotsrgthdLiu94PdIDhiYUllXZVLvAPW+lGRna7l328hrqFy
yX2dhJ6W1/tUkLX1oZjlGFg5Ie6dYItAj+s6yi781ag3PvI+sOF/72Kzz1BOtssDZSp/1WNIyHgw
xJkjZk2HP741X3aWImbL9evPhBk3of6J+sKKqA1fH+ckKLdCO+oDVFXi94Ch8d/BInrpk94VaQH5
+xlIo9vLdsKkop19dyyv90wVcwz36jS+8zQ3nATzX+NVAf08BgmJ3vF0/Wh15qeA2JinoUvCeZJR
5/s/atpLyqgB+j5V7TQsp8hQxQHna2yZ2xrCK4ctgfsWY1CEBDPGYyLKYWq4T1BeUyWUvu5wIUah
l4vu1ph/vUG438plPfLmQC3vpUGCgc3r3siDGImJD3Xy0ONM2yNginwjRrBokhCXFqmL93BwDpPe
8M2QoMR+aqeGI/rqYVG2forFrdrWhd9lUTGe6oW0Ja6F174Dr6nga/2XBYZwLs6jTDo8Ku5cfHPe
15mYc95mGpqnrpFIJivOuMHEgQ5y8x9u+UPohfDvWRgPCgAHs/qamIRpAoZ0BZb+uutf1VAhkSNL
PoMHPxIKpyoMwCG/KzYemjafJA+8fFAHZpmecxJtQRBhtRg8RjrRDXYRbJe5qosGL3VG2Qlm4gYw
WXVKF+HBD0BXiagH2Grjb2tryWgHll9aFtsobfgmcZ/6E6acNMjg0q540ewaxDOTcV55e0qzpSd3
pzyPgocsVclQgS6q6kMjlDYlJwXIDfs1vDXZlALtb+1KJRULgDqd9nHO1Gj756hjMybdb4REFg0o
eYNH7PLVxepFQqAc2JggLYssjAO0ECyjMmcoc7EEoheduL8N1DvMK0zPSmlAlrDDpcJw9dMx8nAd
oFBwKA==
`protect end_protected
