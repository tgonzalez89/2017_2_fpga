-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
pdO6uKdX5szJCL2Q2ZtupfaBYzzW+hviIHTO5Wk0BTAojKLjCmgnKFHv/9kRbDIR999gaYeC4/lD
Ejtq61Kt83FsOLMJWbCvbZd3gMLAsjy4wawsjoKdqF39LURVKwVYZe8XWYn94WO8nI/6gw/R1Xys
1uksEbPkjLGMll0XZ3+wu7npaHlOGHlCDjiP0gYDcNOx5ZAF3reWt4yNcJSgv1Ua7NkGMTL8Js82
Nl0d9ofH8Ydk3TXuTdHrn7wisCYG+PElfyFWctiup9X1oWcS6StZBWVrvqhAImtLDfdhVOe6JdVt
W9QxWJcyO7Fe03VN2X6jCSXD1vmGU5Fd2rgdxA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 25280)
`protect data_block
bFib+jRjBhMqNlkPnb8SWndRdSe/WEF58MgKY7Q5ZmYkn1Lux1u0W7khVLDlTuBZtJ6bFUFPT3Wm
N7lDQyB6+5iGIGPw4l2h52tbniilqP7Zz+NMS7t3amOA37aaIOVBZiqeHkflLKteBj/IRwNKMXdj
9Wm9IRKedRP8ADVOSMFF/StL1HDjzIi1vOHWLom5+xc4BfylTnxBBPEUq959CgduZ7fn1p2YNgJi
FzSuvphe6qcaGH71t3n2WY+C/DI0/m8iwinpLQcrumPRrm/iqhueg8yYdN7BKhICa8BhyGB7+/52
QqobP9Xj5B7QUw/BS+2XGrFeF3LDhmFkWm7/mazif7GpQ8w7P0ra3q4Bi1bCyF6z13YR++e6gbMw
RUGEprrWFiDLZIJM+bZKDAOCMQSeWGxPeKCADvtjbmNoAp89/InY+O0KeIO6iL9N/0+WzqYITzKo
WIXZvPNeOVTZgmX/WmMWHNGhcriRoIQC89aEkjRsLR7ftwwI4mS+S+9WJonMe5LqT4q7HLUgjTc9
/UFEtyXCfay6jJ+JbftrpGd3excaGv8AAuPD1OtPJvs+etdtRgCO1p5dkA+vtLJzIKdEkQtr7kKW
12AXZXOSP7drTgCJahnWY3hcNQzcuDyB6LV72rVZMqny148aSR3mdm4tv8pE7CJYg+nKWc5LaSrV
F0nwC9ETgmsvK5yMcOZ3Zexej819WJ2NbUXmeQOuDjX9rcbMfm7Y5Hr21xBML8ueST7CHtLv3u1Q
7fsdJgW6XqeyczAhbxD8IvkpPP5d0RU/8urQVzEYGHVmMA1OYyAQsblCMgbDjWgOIURo+Osyh6NA
96lBvUrOm5mSphrRCAmVaP7Cp3ND3zUYqwuHV+4EV/GJMAIS8VQeqn9k00+FuH0P5ENcPTVLVNtd
LDecSP2VUpx1tAEI0re5sbljQ47COvO0VHbgXsfpXxumjoZZnlAxM2lwEJPqGNQm/O4vRx+KHVh2
evWrvVoHXeyMD7xUEQ5tprHsv2MS49UctIWXkyPj00L0JDUmjiDA3kPIgLLCBtco8su+D6Ril8F7
UknU2mQIu5iTZIzOg2iJBdYtKkQW/JTG2bfQE8Wz39xBbDqBr4NTgDM6TsZvzTJlXi+MsCFui0Vt
l0NpRZJKBW3+Z0uQlp+tfnM/d4lFVg2NE1rn7mqqzM9MFfxyBoYXEB8fSNSoJPk3NHCV1LGm18Cm
FyCgCXgWjQRjEfAl1Zaea7ABHZzYS6fvhqZeW1psqdb9wsWksjbFUvxZv+6HVVIydojrZfG/lKlv
bdD345y4OQYFvn6iLQ8CA+2NXLbqSemiwchZ0wy0ACuLxHn7uGQXEo0r1D7ax7I9klmjPMEWP4C6
Nf+VR4tl/MTGfbpxxualta0lmsNS7UIZGUk6IZRXq+jWmg8x0Gj2CIk78geo/PTiKZpXlhOQ6eZj
P/z2Hj3NCx/ASv7ZJFju+ryjQydsjKE0jzFk844+aZBJv2QPDeMjtDO+SgrIdOW0PauYPPbHMue0
UFvbSQPYz5ZeI/sO3rnIZD1YnGHz7ZLMqWg9wXJT3IHD/lCyqOunbhVKLSgX7jTrlSBnbCuHzJnF
sRodb7dw0pFUztRLfcbyZgNLTZY8xNo3Rkcp9hDU0Zah1RWzngJrfbesteONqzh67f7MgV/0GIS/
o8o3aT/1mgnxvnvCIZq1cz1Pt0EnLGKVVoRBMPIxyiAZ6RGHGvdDB4dEwnYA4NJXGw1b0x97KPsy
v7af0Yl7P0wv+dWXr/0bsf0D0thZrP+7OZw74XRjT2t+uQ0Gh75eQZHq3m8Hj3HfEPtfko/MqT3s
1OfOecsuKwVNA/etWgm9o5DHMuXzE5DEX3TOuc5whjwVHHgzn57/TUXYtEHt4RPuDUSKYO5/OuSr
8JGHlnGrp6nfp9ccD3XWnsaBBG3Da4tIQsgp5Lax/HGvxWrBLX31AVBBdd/Ic9T2yI+CS7fkqydk
sHr3GmOpJZX4VzFPvIttJxRzQpSKrcJI70ijuJPmLkVWo1PkW6dtHzfLIxms5Fqlinky1pA8Uxjp
+BQneKrak3loRqYmIl0Z3nNgKzn6gjajwreQCBUB+hN+aefxefH8nZct+gPjCDxfFC20MXzvMfrN
jGyqrigDm/bgMuUAbAvEvI1TmDfWHWXx8h68WQwYqnBdbZOySe+Ca8/zvyNzYgwM6DFOpa5HV/Wi
PYoaxbKgr0Dcbot8WKIDzlvn8F7DeXeCgh5tULFPvIh8vJR7DO7gVd0fTuWjvu+t6r2kArXwXysR
WCs4pWTCmbP0EGx24KrKcMjQ0zyMfTBzeyw7JSfiIOyXIFDujqTH6PYJ973Dc/x7o40CzIW7DQzG
2QjPmZna3EiNDl2ofuf1FP5P8WJLqciPTupU/K/OU967u8VHc0HNP4R8fp7z+mM6DaWg5tGc9P+E
/fN8W471LqscGtAm4Q3DIwnxi9XjVGV3gHXFAaCXjdNA43i8/sHWLwSiZaOhUB8mAvLYLKj7yzTA
lYWu0kkd8F/CVKBzHK26cHY4B02KJs7fQylnCpy/hT9cqTo0/X7LFFeNPgfUuFjO6MBSeQ8V7E9J
jyRF2+2wGKGbWCyN5h4AQb9AiycDvd52zOINetMOhhDhsdYWRN3k0+cflzFi6Cua5SZtN0Y5VOUR
9JJeDEEY5U9HDkLFGB7nEk9/Vy3Xh5ELd59YaCpFAOfT7whACdJmlz4RTX32yaHyq12VkDLMXVfK
OI+YTs0AJ+9eSLX29mi8nG8A8t7R/nXVy2ZPNRXhnYfVFpcodn7PKZX+z8mn3ZfY2aGIIQ+aTeDv
voj9IJhnHBne9K6XzLyD+AjfPq4BQ12qEN11rFlQ/oq1iX0h+aNEN+euvXVGbDQiulYz1ckd2XY3
+ptPxIxRwPBmjbKf3qwHq/5QJzmDCm/3oV7UyAiN5TY/hbjEVQWLbY9j0OTtZjKKX0H3tQp+kQJM
sOMJvPFR7EhqS3nfuYr7T06P1gaX9gv9a5B6J7DtfXbgJfaaAMigOb86wvK3SHxNMiByfMUBcS2t
lavvyCJnLOxXCDAuOJGEdIar/zFaX778mg9fTN26BtAg3+jfyY6JprUEEM6VqNLG/5nWbBL/RowZ
PIvHKo4K0ky8+q3/dyVgGEzBhJKXES5dVQVd7mufY4rMjb22k5Y360RlIXaCGa9A80MIFpT4Su+g
B5t+sMb8JbNz7SuS9w9xOJ1fEAAktVU9vwiGLwdo2+8UpDXZYumHvqogsINlzHPnti7c452QGzti
KZsYpziYcKEKJJpPI+1pNWq+ubhPgnzW+6e5FlI6J4CVb61ndD4313gVkv8vuoz5QXbdzPOfKkdG
r2PniipcFyrkpTZsfbWuV4UYe6VU5bSdP++elX2p1rUJNBCA9cGrHViKFsp4kE0TeG2SN0wOJUXi
mzjVvxQpTukwqxdeo90cGXE+7v51freHG0dDoTtTBWGYImwlkJxMygzmcrxZt8f05aX2PRAARoXI
G9WPnECxbDJ8YQv3jyH9ZdeYKUx0r4b4aJdweNhSq/Y1Citz40aTgBfmBXK+5tEgucYcS3OHfVzG
JsXChCnaWzVd/eYRYG+Y5nkdNqXJw5RGR9+w3ZyUmGFWSOPsH3wxu9e32wHltHzbeK8Vvdru8/MT
tg8e9uw+4I5hITdRI/Ms8It9+ZnS0hQu/Kyq12D/0T+gqus76+BgwEYN7uFwS/anQrh5QjVVLrSb
T/ew2oLWjqRSGze9kMHNS2iOJRfqTs+2iHc8nSVGtKANNcu08+e2272Pdi9RXwt7NjaSTIHwfGNA
8BMgvjVLP5SPhXdmMm7s7W+CnXJhtFWuDsucpPgiclTHkozwpqhGBcdgLx0OQnWmzY6l+u0dunGE
8PUOQe/4nQCtGKGCv7jjK/ZrKK5yfdCNf3774vgBGhF0d0j4t2ME9WTj4utcsWqFevrEt0oOFgNT
/94wh2w80Kwqz/FxaveyS4N/IfYKAvaUigSRQfoy4arYymabfBu6rSKZcwtGTet9wPT+Svh4weyt
ZA5c9MaRAWqChvZMEmRd38mkM38es1Ek8lgB1oGHoO0+lXIsg8KapSGUIVQQvkTVw4lEbboedVA+
Mujv5lfX0Qpkv1TzxW/Kr6/I8Lfe0VtWhSTbNtTaCQkzvUT3gPmAFv9/owC8jQbcoRaVP+SHMQ0n
JQFBBL7CTWG94TTCpAtw7Y/feoQwAummCkK+BtMwac1oxfAtmelJKMVcnwFF8ln2duBWtytyzNET
CJ8eR/KuPQGgNKhUmeeEsqLtSVhqs6w/7K83mRJ6BZe3psPwuYPcNn2ThdyXdQYM/KjdL2yO+czk
yPZ3EZdC3tTXuJCHM3Z2n0YNSoTo4wKjEBIefq9d/p+WMTGmK6EdcgutAQT309FNs0h2l1QI3aYh
LR6MLgnUtztyZhfgT5eW7YfuUa91uCwQw8X0blFeGSzI6CnkBlQP171g4xv/UrKYZn8VJ/puOyIu
L5WYNUt1WeLYze7TM3OeUX71Ba48l38ev2NuOYtt02b+j8EhFd19CHtjusbV9hOdELI4oqCR33bR
KHCft9ferH0tVX5aiR7sc/mkVaqbKyCqrclMoy6IJEkuk7DKNi5n51UipRJQtNaTSmN1OQ1vez3J
WeCM5QozXWCqZNHQ5VmadHI8geQB+zBUCRIoxiTJfld2BPoWGzLgSUWJkOy7ZAOw1WGe01qApd9D
U+bZbcBf+tSXFfWfA4tBVnqksEx7DA3EACjbLEKYrLowRZDWBMFjWiBl0goqO3oyHk+mU8aIwl/0
RxpujP5UcHRsludurpXn8TvivLYQYZJXBKQpUViWyl37P5jmyMhrjti4/wkjVJqtZhAwbTjK0h1v
yg16owZE2FpMxBEV84UfsfM19DDS+G7NEnYl5mg6FdAx23i6xkqoOCphechGjoRpS/uHzfMOOtou
NcVnkP9zJ2SfNBKhGc2ByC9gJ6zLgt62ltiZUwyL26BGt6BzHFfqcHidHa5ePe2HQqNJ1pWHMnS2
W7BS0lEB85GU08dYUm5lKP3gWoiTNy8a0CrMBCk8wpBAmgiywrR6MxEmloiSCbGfXqwg9lZKL0Cm
Nc26sm7qjpp/c4yWxJ3QtvxF/QCm8V+sSdqIJgw/NFfwqHlhwBmO9ALatue1+S8rchRIDLW8vILM
qz2Z0mMS0KIH+alA45dzN22qvQKS2JB/TqLvjc1SM7SwZjj0jy/7o01JLroLW0C8UnAU7laPcAlZ
EHwdqkNDdX2hdLvioOChpX/RZnZk3hDB5O5sd22etdC4lMvXdL4gctj+1jZE4mlQImPXi9PTCTtP
+G/4h7tSIRxwPtvPayrJFD3sSuM4ccC9ajVqrlueB0kpPxPTP/kMgpxFaCspRbB5NkHD3481AKno
Yh6qXOtQTkGK76JmrW/e5J8Wjvh4sJYepiOKK5z5P2Od/I98fA7kfHgbFx7dyQtgPSmo9+1zUsn7
KzQu7ttu5qsGGgMb0BcJy3q76pdohtxSviTV/cvWIc/HW5f+S0RebfUSscXYZqzL2PXMgI8jDrCx
RoHhnZn788lBgL6A1W2F8LwxH2IV+JpQp/rMQMJdVtTpTdpg54XAZ009Ooersq21hpSR+ohzBvUm
+Qut5B/sSsIfIQL2zRJlT04D1W5ODGsrr4bVnx2L5igfQX42IEvA/JJDEfDIZOpkiQiB1cGq6Ny2
ZJx+5f6jgy+QsJZSDEINHX7fXe4iEaawMiZq4iQQgMGyRwRQ3nmnlZxC1jqGrycZwSNc5ybSCMM2
9rz9VvNyh1K0rNMASxaYGjJGpUzIgWNUbZN3CPCZJG5FJZZDtcWxyhgMf0iJXrNUnCp06+nXfPyF
axpvew6tYzBvcfot9EbZxldaHaS/iaV2rgqkngGU6Q/6LADstVnsjvRoqYytUXchOylZUCrEbmL1
PwLFmSV1X9oaMeODgYkfeaqTy3R1DYFOc3TdnD5Xsdy1vE0PzqJihmtROnj7RAakMoJbeGYTYcKT
datfq88oKicGmYZwSCMh/gDKG7YJUWgv/6qnTWmeowyR8LRHYfj+3qF1GusH0vpg3tE9SIEhvMSw
gKek7FPJABLV2OF436LTeRfRWT8jCWXjmxSgNObm3JVE04ERFM/xBK9LkYfIxOdcJ/FhWbGGSxT8
XpE6onNXPlBcTLm7J6Qp6lVTk4dau/kZcgQfwAHm+UYhzC2tfWdPCxln1mAUYVPGJJBBP3d7XNOu
Ltb9C21k+ZlChcrOh1+DSC0XgFGBrv7RwFKd826U6rJnjWW/ai2QyQhrEsw433Dm8KxzsP+syMmw
meq6018Bb5r6mKQk+U+f153Du754HRp1pQvFXkRIx9aAl1jdPNVo9zfJIgBfmT8YFGvpHtqA4mxZ
XmPVODbg/irp6LjShz6Z+E/V5g+ml3tyjcKeF/ZLJj1ypxh4KXQBoDW/zTLbx4J1tS6jAKQPCrXj
UHgciF1z7Z4365gCQSFA/LeMyNSKNsTK5kzKUie3d4fNJlnv6x5Xxr2NlcDXKStiMFVAxVfPb+T7
3nuExNqtZVai3tkIFNw+PLLCiDa0dZm6VlsNEB7Jz5J8CGAmBKtF/G+krEeqfapHRhBHDOZxsUj6
CZcY8f3fpqC5s/AJW/RIkg/FW2043fBBapIa4TePKSmT8AOa3M269OvGBcVzgitMDrCVDKhEgzTF
Ikl79h3wpOwQCWEmdDOnXxtOB7xmrWjZ5qRPk8AddbFltCCP32AeyVB89Bo8OZptrJrz5TdIql9W
T+Hkt3RgKNAImSfwY2dwnV0nqOTFLmaZChW9JrZ3XMcBLcnxqKKaOlMx0oTs/iSBVIsclGoOUwCl
v+yD3P4KUyZHzvG0/mAPlpEuJErPNCSCj/0p9qB87ekblwr+S0w+zKhr/9ot9t6sa7zf89FHuM4r
/PGaHUlikyRbVca+EleuHtQ20RwFbZTULueu8+RCB/Rsh9ndM5DeoRLqWw4TVH0dI5Lf6aeZ0K1X
Jv0gojzzzNax6xZbc3xirRtfAZOIxraPYoJ4I2Go+mDf29HWYTmtdY+kdMSM+mH3IYE9u8HZcSVd
pJx/CksqYYiw0vb+cqGmZU0719TS8m+HnkO3S5N7MNW1VwgE8Rs1+lmlS3FEcZcoLQN6kNkhNuiG
Lu7iVMNorBEMcNwC7Bavn1lKEkwxLeET5VFNAm5OLNEPfO8VqqKCIqmJd48lPSfcz1wsHQkBuOyp
UrMQvHM3klVs/38Vw8qDjBF6lZtoABOplKBfZha+QSNAtNTNb/29tYYbM/zSNuLUxV7Yk83HGI7i
sbOyFCKuFWAJXHeO4l1ETS388cqqeUwivHosph2GQJOPBi6LDbaJP3bfX9+tX3b2fF3WTh98c9AU
P6hXPkdddUls5xlBE/RGU/YSg9X4gleYSZ6k7DGhWGfAwOf8/KsAUEBCdGLRJC4dDp1a5TDsS8hs
4LdTDEfsIwcL3IJOStgmdNgEIHMkF7PjBUeRa9fkQpMXjl9IO/qE9mAYxuWa0P/TFLZGq30Fuy29
Kv6My1YnGAGmKz9IemddL89kHuPefSqjaIuSJD6Y5Esg1j90fOlKuhQ7aMuR8etBoS4tYZ3pWDW3
TqKO/PRfbqaLuscyX0CkeXSfQlzlcaUdmEEVzdPeVkI2xxLIGONJJpYdOqpohcgprNcfa/qqWiyz
cqeHnXm+0KwsplcQ1v6rvrb9o/1qD6BI3XXqNPR8z30H2FLx4C5G2mDC4SLOETiIr38VLSOr9Dbv
J8L8ypyaUKvPB4M4F6Zuv6KRkWVcFPbnaJ0E1/LkQJwb1CJIjd7SDqeaHXmUe/f925PkAOG4Vsmj
7v5NvY/few2rubiKs3jqb09+7RVCHfBCtA7i4HDGZtHoUsOxxsp2lpFFOOT7k3eyl+wcHcLs6GvH
Pq6lFZE2aPQp4baGchFf++hA05iUqxKV5T+hXYvFrPPQlOgGwZsyZ2MUP1S/OB89kgRDkwa5Dt//
Yc3EEphA9Ey8DWldsUz5DWkPL2k8U0wCnHiVws5Moa7LwEAf9gNpvocpJt9AG4GAQ7MkGvcdhJnL
K1P3zh7DKT5JNo5aeLGCWNkVU9GuBsIs6IYxYCttqO8+mKW3fd7XOeobNuMA+usgnQ1qSH7Q4gQb
owUDsvyegUuTL512ej6V3rBVmNIhRz4MbdXxib3FCirBRlcLT0j46FJQXld2b/xlj46y5LzcvxdE
4vegcedthRgPLtC+7CDySFB/aYoWqsAjyS+TRH3xIMRmUmjJq2zMkRRODaQGsGvS1Gd2S54N5nOf
0IvNKPbsunNfftdGsPlLzPg3kLBULOvV65CXX9/QkhNLnc7BCR4xs6u3reD8jL8sHbzahlw5E5yY
rb/JiX6CFFvdNkNsvAPhlBhal0i6fvBlYiGWYKvZ2YvPvexUV4tIIw2MPy16X7AlY5NytQXEJ74G
t2pSrKJ/YP1EkmqA6bsG26i63r1wV1miLE0dQYSf7WPIRWXu/NNL5aFZmgEFcpvPlc3i2O4doYcz
+tLD/TOPtm5OxfkznHoe01+JSbIJ74uZCDrziOlBLiy9qMh8wcXpQe5c/90Ckgfg9aHuUT4AfHvf
fwQyftPmRcrIMtr10eURZhweNCK9jT2TJtX9UX9rsUvgySCG2iq33UstUv2Ax709CtTuObV/VYIB
bHbT5YqN9tR6wBs/bdtuum4tADQPQIImS+68rdpLw0p3PxBp4av+vC/MxLwycrkO/DbNxYCqvORW
/2eJTf71WijCje886XL+yspZE4ernrnKdeCwXe1ufLCiAqCfz/ZOUkBZq0ihlWO4eS1OgjW9MdWk
oLEr8dxAhFcFeBms8anSjUcyQTh0iVahSs+hQDHMMam8vHFi8ftx/0UqspckoDqTLO3CSWilzzwH
jTGYWU3FUOn2ESL2kyCnTIOlHUpvK3pdRteVIJtO5YBam+wMSYg5KBTqGrGXoBL4rRMJLHZ+MzQm
kO6gWvGEQkJlT2B4bbzc1z8+9sY5N2N8feeHq9r9x5gZhtSmEnT1niHzatjqOFuyIxrKbIJKjoVR
NaE2Pg+LXMSYT+iV+6fQPKtnn9CxqazwcLGCN+frlOZEr5NDxHgIn6vNBhaZj1iymN7UeHjV7frs
BfgTGeAQJPny8kpQM4YNatyq8DpDMTEr01MS90eCZVegIwpYmF4FfPMG5W/2Kw5PlT4L0zcQMkhq
xJl3oLrA2NtzH8zUi9WsHMtamk8L04VHFFWIw7ddyDuvNt/MFAb3epmDDXYUzQmUH5sjdIvvBXRm
NWJDDfUsGK0se8RLjzv1S/QVFgIejvIqc2h1t6SmjJHr17Berfh1R9vctIsQ5ul6JujqtewSlEVB
EtghW2NraAdi9uC71rriClInr+wkj52WgdVJ3TLK4kggzpf4dVH2LPQKql1qD0w/3GRNkHkd81Rn
afOSffOuHdvJ81VE+18Dy/ThLJBUGh8ckTD4TCvKLnrfzhHRp8Cc4ThQ5efg9tojMH3lvzaP/vhH
1CuNo7sAgQxN47u/h5ZbZxyLn0mMCdKMBz75335t5jYHAqeYByg6mVJwRcDhX+dZVJ8Q9utp4qEh
r+O9eD8ejK1XNgSeTfxFVEzRMt4B+yg7NCS2dcha9cNGO+ek2VniEGGUQs+3kiSfezp66c7lsBK8
p3yIs1Hu0VE1o9zcPCNwNl1GaC4hcpnRO9h3JsaKGWjkP8W53oo0MwsomVtY2tCNk46KgzW5RZ1l
yFRnG8HShgQl68eaeQJA0Zo5U4hvpfLdMj7Fqq7XUyZVod4Yjx+6JWbKwg4+w8/8iKZVKEZ0Nu9q
8Gld2xto0Kpf3d3bLDMCBDdyWtInb4MnN59VD0jjFFsfApzikC2fTI/9XM+mjB/LHNu1a5fl0t6X
jY/OqlcHV1oi4jfcTiBkX0y8mp40jNoFb+tt6MonaEmKJrfdfGbHT00I0qagKCqTDSi4fvUGtscI
h5tEsPZOcIKHVbYXND7BuME9EzzGo2xC3URn6pfvV4es9g2rG3DVxET3Yb1Fmyje0x5GxUjf4C3Q
DNiDFeaNy4mT/hPrnYR5rULtLiQgYXLSoxzSG6WOSaPm5BQmuverx3TEYi4J8T2APSPfD90WfYQx
BplIGjL/wXv0jagqV5nJMR3pgECs5cBRnh51MbxZlKfI3XIcjvbUTY8nBVBY3Bzjh+pogRQ4wNhS
KFUONqrO8jvWVF2vUf9SOscl9f3FnzUDV9s3+RM0xR8kn2RIHE8RVSM5cPCAvjgvVLAhdoonk0qE
N9PlNQBbtAnF76htENp8L7z7ZBsMtd+V3ISMLqLsXVW1Hjw6R+gHxKqepNvvS1Ew1PZAcEpZt3l1
ba5q3MD9/WfiG4sXrGdIyXIlCesTWy9/Dbap8YYAkkSZHS7Q0dkT7SPvi39KUtmJd3Sddxnntdfb
DZ0C/mLYlRzgWcYkuY8Ceo8xlS8GTEunbeidgHh3ozzJi8lB4NWmv7HZzvMWZB2K5QID0tL5rlua
Ay1pp/s7jZMfwyi116NVnVxfSkn7H4ra7Ght155qDw+K2jxaN2glmRyIo3XsRfybGZnSBAY0Q/bg
y5hp3FU8fJh+W4QZYKwINRrUCmCB6cNEMjhjf98lLQ8EO7Y+QyEx112tgXY9x1/f+bUgYKR+pIgy
Q2TC2axur0JIbHwEBGEkidlJzAJ9nsqoixo3xwATLk3e8lsXzm69xjVuxvHQVREo1zC7KnQ7DMsh
ZaZbsOIO5Ami639RHSnb3szhh1JDkB6QJMq6d/e6EcbV05mXfBNXyQdY83A5C709phoJrwJhoNKv
tstNe/1i3gpeCo/Vw4IfX5R5xDB7HOjmzSXyGUlj2csyjbr9/bJXYPStcGOKJjL/AXmabEhVBtol
8Jd/D9OgvgCXKRmUeT7YSPayfvpiPoS3cO4NzErsgTw6NOl6YEZ6044tPBSjnEzFkSyVeHdOQa/u
8MXzl6UXk5T1sRp4+C4qNPaXEB53LmL7tsyPngaEalMyqLlHj/2T6t5oOpzGb1wWkgdVOldelTSq
howeBxYECI4RTdFCGE+ZWgNanIkzgIMplGtx9W/kt8/xifqlO2vXYO7WdFlP/qBWHFuJeXH7UqEu
UAvqmQJRzTvyu7zsyuKB3GoIKZ3e0tIv+ipSLQqZVArATysA+lbWrqKlUvISqjfDemZsayBo5LS2
NM5zeN5TfZxfwN6+JkbPjiaQWMV3KoD0s3PHFJXrJ8eidCQ09j8kxMz+fMOXJRiyASeHvfsZve7c
lFsD6j8GPvAyaA6xr/xhQDRtuBUNvOmnndWH5J8ftcA18se5Xku0moOvZEgNGs0oJ2kk8D2JNH74
4ZGFibL+/qeyQreoQFAay6B8Y0prK67gKfVjl9TSepdg7eXeG+nJI4PxU2c8D67fzCvSyW1Vunm9
Z3YYZAOWFwNkVbsI4+vJkqcS6yR98WCnm0UJx3mizyRudYyagoWCe/wheHttPOZmZ+++eC2Wy8L5
xDHAumWEMbOyYYWOXWdESkaN/kvXF79wa8zNn89LwMXrWhRv+RDpuDi8fheROzWRp5icavHiXMkV
nQteXJg1X3xN1loiIy+s9new2vwuZXYhDg2R39j8NrXxfz8QfW8uSy0K5zhzxycfzE7tJ5RBODdF
uj/XnhWfzD63u1Q1Kw34y3VhTCo3EXqctxi06IEFcocgbU/6oBR8nyaSjAdOLuXnVKOHhDJDcukh
odChnwCPER0JATBDjh3k8vfhQgaCnqS2i3wMLVw39xugi7H8GRIw/YHugLn6YpOd6xcTj9G1CG84
mSxpZqoQqoOqGwAXAgYmuuluHib3sGTpHUjXq+E1SEkoAahlssTbOjPpibX5y3jq8u6XZTJvianQ
yjwkFwtyBoa2+jY6IaOKiJHrxh/R05RTyDMeUlLQ/G+izc+o1yM2ykVY3nbBrXs2Lhyeeq05Oez/
DZlYQUMUNJKT6i+2HWDVhqc7AKGYZw3aKsVPkCm1bQ/owK2OkzTiswai3wAsA5iURU9JtEECgwHk
HIIDBsCqpMBYed8mFvxtwqZn8+hT5daoz+v5XgkNzK2uKbdv61eY65zeXmn81Rf91c7ApewTPos4
6M+QP4wdF1xs2OPn+DdDBlD/F2jP+sBI4vYU6NKxVMklXDyvVGY5YOSY0V9Q3EIqifA8O0/1tVr/
ThlAlK8X3B4bSPmrhHtz97a09Dc5C4icjUeYFJ1gb5nxDGJxcwH5lwiVvrfSEdnzHxehhpGMGJmm
B3LXurCB8pndaq+/Ao+mxoA5K/6/ImsXCLrXrbtzo3UOl4NByDmRGg/KbRI238RedfJ/EfHj+ED8
OszFKcrT/UZofyoRqT8+luXoOEEYjGovNsW40XPgIDE4/yVd5dB/f7g96Y/ant07O/cWgHUdT2mz
AxTMoePr/YmtfI4UNGR0PCWPg756+b/uXW/fRRhfjaaM3LtcmVZ6ZcRLVnUN5tyPIsa93+uytqSF
VLPdcxnJk0uhI9vNB+oXM5z2kRgulCmF/Wy579Aj5vFH/LVl5oHQGR+MDQNfe55iPKywihJLvF1R
CsHfUS1l7VYOo1hAFJ7MrTLCZyNc8IsB2GjCSfgxEdrMzDAlvJ8MAcaeeBwTv9QYmDKZq0nVkxFh
VFXaqGGJmnLV8a4UOMZfDBptBuakkK4HPv+VzfPp26O4Yvo4u2fP3wxxzbfTTprepUeMM/vDxrW7
HItp2VJiXLTcS3Rucv8zvBGeJ3RoLRYX98Y+pw9g/Gch6+8SU5ibNA1PazOdhnq/6NvQdli7R2IN
gjSFGaaDSq09QgGp112WHF05u+YHNhhlGISp3BIAKTQUNKxT6j+v7hgviF9AOHuG6dnytH+fL7qy
AM7a0YPq/Q6x82cU8pXJTVXjJfkJk5suUJzJLjn3AaXQHyi9DS5sFZwrVfz3tpWw+AVqL2WUWDQH
Y9KoVCVbGDG5dyTic5pZF1ms7v13xTOvck2ZhyW4E/p20oF1gTF4Dlu9oMn6iyecx1OrdAhOp/YN
YlpL4CgYaH/rBDOhLw8RgBiZnx3YaBY+HPrYgVYkKD0l9Hn9U1yanIBw4reHdZ4eOgWXLB73GaUM
5tU20SA5QUeBvMB4aTuiWMOmcIamxRqs0wPcKtS1raGKfymPN7FJiJk1MojRY01W5clYWg6jfcTx
d5SUxBIVcpznICazlzHpEuH8LZTss6aKsjYA9LQTkuUxrFIDHOjI2EDzSxFjD/xRUrW8WJaHYqti
GxiEeDjXun+gdfgonjfI5SQHT1l+k0sSE2EvbK832kNFiyj9kJ2kdBa3xiO60O3E89vgNok4MZQZ
yHQ96UGaKnm/a0+X6B6F0BaZnLJPU5qbjXr7Zm0AdWo7Lzcbt0aERku8RpWzQS9yCzZ0C5JLqzMz
du4BNx9TH8k8W6JQT0AYqwrt7luOq7idEPxyAmGn7OFM7no0v14kt3f+euW6Nx82QZ2FFTTNN7gk
6YEEdZg4BRuoig9m65qi9ZjELAm75bbsv2GcRdQIcUVri2oVegPr02Z6TdJu+B9XmXno/e8b4iaM
ZgNLt0rysNgnW6nRniHKfVc1Uk/j0vcHT1kKLARkhS4sodO7MczZwegEn6ngL+rWBes+kakquy+t
yY44h+Zi9NwsaO7NbsOj8R75JB2jCrpRZuXfS8aA881wjnnLSn5LmokC8PN1xNCExgFDXBB+i5bp
XTfj5sPtfRU4ZXuYDiCfsg6SfDFq4bs2WuZxjLnjbvUdzkCIL5WR3wkJ0cdO1V+rsyNoj2LQf0hu
P8HrPtEdoupMTHriWisz7qPkhe9IatHKbeDV2ONdE4dAhrkH7Te83/7QKD5XxObWnuXluYPzdCiq
/nART8YSaZM1eJvZH8cW3qhyMBRH0dN1qj/34Y4CbM3EM8/daJz0oQoG/apP6DV8biwimSdmm/n6
BKj/1x8NnxiqtlM7UQYvf8S1BBk1ykOqrOsByWf+96hR1lhgb8TMaJX7DtkP/g3Iw5cgabbgpC75
QF6/Iw7CTeet5ONeBlnxwf497k+la28RrMoVRn4gvxFnU/YYKYrG88OWY/lY6V/8Qp62vQPCdaZp
o1G1gNm/LIgoemoGdbEhZDQnZUtf+eX6KGDnVwNAk4GpMV3BnTgXTe9xQ7st/zeYzSj43tZ96+si
9WezpoG+3mGDf4Kek3/rzSNNdF44AgUz2MbX1cwdBUEejXDyRv48zr/ksGRuPNr37miozMKWe6Uj
sDlJhc8rF7rQNLS/676mWE2nPeB0FJ0ILZtNosAgldXyuqep3gCTOTvbGibg07e5mqFspqrR3Jld
sKyi62m6U0ZXSUwc/5grJdsT92pE4bnzN4rMB45fQrs5d+tB8pU4GoWUSDOSDbWU2kb/UBn+dERi
6ibU3rtGGMn70Ti77+jLtQnZ1fEznXsmoVHNzoYTtkC2lY4UppSmmvDKgtc+ml15uOaslZf1EZ9o
gmp4YBlFLky6AaG1O7mC+OqGMapHHNNY3wPUGTwH72pRtsPCI3TUtPXJLl2VYH5rsgkImJAgVLO+
iOWVwwcjXsj7QpUIFQ7oNsTMTV6b96s2eT9u+AMMdWqPqOOOw3dm19UVL83XY1kbrFnrZPlDvsHi
QjQfdHAXHwU7MBjyL+G9dOBBXThPs1BhOn4M/7hNJ9bsc6eKRkTOzywdYzkV27bxPwHKCo9fSHyr
8UFl/F+cFG935Wi8xp2E2T8mk1q/LmEFgo1Kw9OiOqRTlUwyGTHL4k8ZUD7J+pQjx9tc7ZQQLEJW
na8CMxFg5vMLRcoywqZc/nHXTkJvE07YKTLiz/HKHQstIZr27Zc7bVvOTL2UxwF/TBr643heMz8w
0NFuqTsUQzx7LhFnKw8jqYIJwo8fdHPddqNh5uRqRduHZim8PxW+knrOU8NNY6+VRGaarMZThEL6
zbHQwcKq5aWWFvMLfJNem7fKmwXtG29K4FtSTthYvGjFcS4nPE6ZCgfWqwCH4rDTlkNIhLSSyX/B
tsVnszyFKaELmu05dz/wEIR5huCO7uDGyR91kfM/GmFPXqED4CTtqP1NsBnPyjU4a0W2V1QiTFcx
ZWY6+9gQufgJpKvErOC7cDuyVXQoMm5wAN9AyFl+vsof1TkNyR2f1mPn9THkcJuHmoMtbSwsGGRZ
Tg1a/WOkc/21AI8EszRhI/PL1habUbuoCYWjxDTyNwiYLJ4tiz+SaDxx/+AVBptbAdH5raeAqfCp
ANXSnCQD4dma9KF3cxugLFo2/g2xU8KmxQHx9Bk2Keyeq6/7luilm2D4nwrqHrQtTf5FFLGlGL+b
UNol380Tugmx+0o7lrPbbDaQBImGn0JR3BMcXWhpL1PnevuLb4B0vPnXdrVeh3BbpjUVVDuIjrsL
VzWPT69rw2WF1C5p6SRjx3mkXDOtw9qL00mIdhcFJzxeR4zsVBc17Fy7TYLs6GzNBpGN17yVTm0u
4EjSMluHFcTFZYVrdkaIsazJyTGl2P2ABCDCCMscLVdzN0Bj0gN2LpB2J6RsO4toZYRqBLiqFfld
YUb65FFB9ryYpduxReskqPUcmZ13bZM8pll7QcVsnNAHD62yImeHhpkhShq7ikOBXa4ZDSIbpT9g
BFmQrl00Dt5CY0YEkUC0d/knZNosvu6x1jXU9NQvxsN5xWiRZjBC7yx2SSwI8eAjXnerGgHqOpRN
9SqyI8cpf6W1czoPP58Xr14s6N6jX8tXMF3PGo4yB4zNTRCp9ex/wf5XYwNf7Ulccc51QJwD9mYn
b/ajiUxov/WVjJ/P8/Y5OQgdtHKVEGpcsNGoeJOsHycFyMyLAHT78J3RLxgteqF1Mj+b40FF+5XT
gK1Qp+tFs9X2ARDyRHfsnkGT8lftSxVNMufRnbepL8VJp5nYAUgcIUVPa/jF7BpEEnuLyDm2glnB
VxQMRgIMd7kzqhjX7uD2cFWzmF3AeQfRLN454fLQYxaoJBVIHUqX9QHntxLQG+IEq7t/xNjNnxIO
OxTYkDLFJ9MX1SXLTF5PbS1qFn1leWNRXHP3PlHGbO1NcjqD0Q/NIpP9JItIna3NOvzplV8OYHHQ
mzCZUizvrwY3cKCpwZsusXMQS+KjRQtpuD7CIrwOLfrkd6eWXSZMkUy6xdVGReocZ09l+lF7VWs9
U+2zz1r5qWp4sM4FDLWAXr2XWVeRJUnzjdffDWbu3B+lTYYa9nH1I/4Dfskt6S0kP9yrRpH/nqA7
FGJPntGFd698M1j1u7RK5OgqWNQM5H4B8ujG0QLzwLryeFH79aEB75/vc4zL1ueitx825oSRZgdf
ly6zqMhHC1IMp2zSH6kcnxdqU/XyAhYdCofBYB1PB5gK/cZ++4RShoWKhLY8N6a4W8bw8Kapz0jm
xg18fMfzphtRpnVt3EZ8LcIdNEtY2p+R0dJwmHQvMwPqDTZoCKsEAUyRcZKMYr2zxjAidN+vkcH3
N8xPBv1yEbI/kkYe6eJmQolJatB8+w80rAdp330JRJHKTGN6ST4TNQXHLNKfLm70VN8CPZwNDxlN
2yB7LaL0ntQsBEwpy2UUo3/cOd4iAl9tI7g5E0onuVRp+7LiiGWTaDaRM79mYcle5AMvjQzaknbr
GfXeVrDbDCGSU39xmm8TwwjykgtW1n798wWSiEUr9qj75lVuvBW1KZU6Ptru70uwnl8/8hR4sG6B
fF2/8OR4Lvuf8q1QjMsdL2TQA0oV3tAN1l9EhG8aYHW2HMWGrbd3b+J+hmihEbRV7JhZSm2gsXk5
4raSzvZ/X5eg44mPJoHjFX71kIdb7JtfsVpJmFMX9SxnEFJtgE64WGus+xQY2I2ysRKafjWPYEi4
Uk4rUHyePUpRGnDhWFS3lXA6fGJC9ybGAmCWaDgsl/c34OD4PaOF9gFh7qwiZ9JcWZXLdfxonHni
xgBG6VdTyKRcPZYDkgFhXTcSwtT/N9gvE/kSgxJO5nyOHQeHNZfgznaq2BThJuhc2Z2s1gbeFzWW
9meTr6f+0IfNWkI0nv1OHHTzXb44HPL9kNqNR161nQkr0nQdiLlw6ab3POvwXSyYKm1sXTt8aD7+
B9fA5rMEd/wknDciJ/ARHNFC4fMoCqcLxmyZ1TzXUB6+5Y8oJB52inQu365ql9f1AwT9g1ZjfO0R
clqAF40zDYLdJMgJPoTrE296hsGOIHoTTVUEcfQEtf5E/S3WFinZ6i032Wx8Sm8hLt1OhVw91DEO
AwSB1X+NIYujsYeRkehXEcyxQFZt7Hc+TSs2RmtvLXRiKnVuu6jxUBf8QiBDYUj79wAP4ABRTxxN
g2FMPBfr08/TGhnz7BicBngVLqDDcr1Rp9XyUPSRxv7Wx+rVvJZ+kVXrz7DKFDr4lQ+V3zYH8NDE
ZtyfMXOVRKH1gSjj4iFn1xEEhWnUE3DU2duLMIx5E8c+6iDwW8t8Be24Vk0xyb9eh6ETFAMPu3Ym
EE2l/AUa2le5r0fnDb9KG5uu7YLbAPUDBVIvA8A/AeHnYyQDkB3GBKYMtHIilArOLMa7Aq82yu8X
4QRxHKhB+zvt9d1aLji8YTJWxcRh0cYdWl+MsqLB6NmYxPFGoJ3MrDcvmc9oQtoqE+V5ueskPAUo
bSOwWaVHxRppiGLCG4RprhQIepQur7SEiX8UbR8sGc8MiZsZmHqiV0zd9SNa+21gG3UocuuN+iRH
+76DLL3eSKhuuycqFEwXMahCYF4FdQNUmzlwSPkCvtNkfaOG+geVJHn4p6feXPiGuCEGplvXk3F1
5+97ZUGO15uDr1qoSb3CNne3St9OnacLeOirTGSlr9uRuBx7w2Pw8/LHEE7qsA1CkJ4aWSj7ci2n
+1ZzQ8rGRLNzNBvs2guKtqOXMbaNokvj7BfQwbzrQ/mhKNac8HnDfpAwp9yCpH9NL+EUAZBTVq67
rE9YlPRhsTdeCfY2+gKld9rC3qjhJ1fqKbQVMereA+Sd1Jnj8DWiP8cb6TCyXcBO/GQ7CPhMGTb8
3U9cFBABQJZtGnA2r0O8k3EYIY8TNptLu6KVNBojr7H772NeKCy81bHKysb6BDHGlGp1/S3/keQs
qVeHakVmNgjj9F76islo9lYLPtgyzmT86JeXOvb5V++6f79l4JHrQBi7Mf102XA+OlOXynBuCIgp
1MVlcIcMUePnVT9n1SmE5XDa25QlZkfQ5ZD8/wQnlDdldcQPwHBkN6+YPTf7GARYTCEyc/iet+sJ
KQUjKTVATJ6/ZgHOFlqz24lCRaQuHW/S9bqZCR68bZIxAjYAKrVZnKJPPulqkVD6r05A2qh+BmZ2
SuFBaucuF+TEL0Nu/93GOK3gOGONw9wqtdJuVCygn9mlm2iGI/+1y+GIPChojF5ug9KA2mRNGAxq
VcKxYwRqwom456oUBcGOKfT1dAliYqF8vQHZlyTolwEhPpx83Yw4WuMUJh3E6mGcPJj6ZDTJTz0B
f922j5e3P5eB9jMnhF4CX4GESnQUx/euN2vPQd886wOWeHJbAfORBd/R+H2YzRO94QgJzEB05PIX
hyi8EDAWOI32pOM44jKQ0ZGykR663eFm/CGDOtWr77mYzBmrV2E+F1lzXy+oAWFC6G7lWIdtSoF9
lSWRPtx9R1dLzkZUiml9hikAJ7aomhbIbU9/BA2Ao5LaKk57fb0ED4OgPp0g37uwMoI6VX9Rq2u1
ohKxwszywAWaA07aQVJ3kpX3eIVSwNDfstv2ErUkHGLofIyPMk6GwBD5VgTKdHmku/RqX04I81kv
VnTe3HR3AvGQ8BMCpgIvp0k/fuIDy9iQrpImPXusRUCB/Q0PpJq10e9XzhWzrDR59H+ivk0z6ogc
e14+g2pM/i4S1FsiZgT1DsN2ZbvVN8hZP8Y5csczDO2W+pek648asNL4QVuuitsQ+eY/c9shmaVq
7jSlmBPGrwy2HZu2Ec7lY0NA2tSX4+1P+R6DGBB9z5oHV/ZYBn9kj+e0QhFOAmHyFOv86MA0fmAL
+ZFETpKUvRHuOrxPeGpCTupQHS+UCftor/HDfR9CzmEeAVyoaDmyUXUtyrAV5grBmTZJV9QkyiFB
SovQJb243WLMd+NBARIrFHhdLmiPDTYB2lAMhgu0RDJ1B7mivgSMwDDK2aG/x8TSNsEaIcnr1Qzx
uBfql5TugNOQ1QE1ZpY3Z0KYJG+S0kCbGEb/2wzONfnxf0WdPS22rxjOJYwDSZQz5z9nkuWRZsiw
uNa58CDO8ASs6I6K1i7i6TlnsJy94Y09dfCqgfT5O8xB2eGm1YicIrm9DaubnB/C3kqNzUeoyKmm
tUBC5a/SjsUCsYdxMIkYkUIZuaM6xKIsjhJBkGuTPjrJJ1HWI8D6Nqdoz+cAdLS+GOMF++8rVzi1
Q8B/DBryoUZGwolaKVB96e4/dVQ8mmeGIZF5ivRKPe/VkbeTGvJcAiC0t2O4EJPyFTIqTbjmgKD9
R4W/LEOXamoPkoeaoATcVhFJyWjcZwE6SMqkAnH4OM8OJwQ2V3ZD0JeBKZhETPat/6dDbRfasvPy
3fRPIWDuBXQoP29vCtJqinUHbFU702YQ6EIEzJXTU0iLDWlLEZTqL2CHjGizPMACWDdYPgdyKgBu
a8HwhWEOqvhEJm6WcjUVSfvCsGLCLUowZ4wFbWS65quorFHWtzX971PB2oCdA+S3x0+4QXkAXtMo
M54l7cILVsiubkxMuJg/bAvtKzy6nfDQKni4pZN7BcAKnYCXOi5NM+UwJW08cX71C2C07GPFSg05
/XAws6xFFg9yRFNVpZaZM3ubeMpd+obBkPbTu77OFpiUJPfR0E/6SzSz6O88dDXdcqJwpgPt4Dxv
/scaMGsUvoNBIFMVw+qND4Gw/kVNAU5ZMegcpld3SEDfAd7nMqtPQrTTXAvbJV3LXUS+Hw++F4mU
8RjlzRtYJfyf8jNC/kXJYghl9OmN9FHesE1/4rj02HrGlqNc/j2HL8IO/kVOfXJeteUMQmF0L4r2
ibbEDDGX7wzqweevHI5snrK2/gbrHqrVHlwuuw9nBGIe+d75t3HaqrL1NBr/uM/SAG3wSDpmo2n9
qZ21i/jr9swt7xvhB+PSdj220Uuep7F9Ie9sIhKP7rrObZm+1IAyFWmpw+7E/x50LbDqxf/uGguV
1yWmRuxqVd7zP2WzgNKuts+9ZN6tkIJ/3QfwzgHLWWaJ0+uyn4IQnbCIBrHNmKSaYZBHTm+L3KU5
L9Ap3wv6m6ANHlM6Yx5xQq/ozwHPS9cRReIJIvjUEOaV2voeEeXGC75IIx/CwJpBMf6VBIDF6qPD
FWyQ5GhQxwbL0MtZVbIZHATYTYX/4uBjaOht8QpPgGtov1JQ4+UDVKB1drM1EnkdIlIX/9vX9cW2
mGlP4kiTnkMipKcf9YPYmOW5vhwKM/Uh8ij7r6hbAfUjAJzBODiOs9m0An9JFeYU8SXEzNqUnzcr
s5oxi6nuDqugl1wQjyakMX/9ErisfSIC5BpcKKy/cPVCx6nsX37W8KejNZEDQXwLFDAYwYONwxFW
18elklx6Cb5vd+hx8m/fzm5uRKQ+PoB2iqBBBRDbZm4KnAulJl+QNMiGtxXgPbi9Ph4FIfyEglre
yKy1Xe8/D5RDcMjWi84zqux7tbZTovou6tULSPirlOpFyrkVNiZ00WyOLAbRumN7qIQDJpg9wu5i
0LJZSLAFVPPjhPy3vOrCLd/ay9kSZkdKy9HiBC3fnCvLeppgFIPE0xpvwFVtK/dPvRK6uWHISlct
T7p1rS20opp6dqFjT3KOn5OAJMMv+ZyBLaJixE42iAMLjor0ktWkwT8MSxDdNKT4rEktgAm0RPKY
+BqsaebsH8NVUBs+4RmkYp6pYWQWSeylN16Hr3rG/xgmKh06UJ9B/MsG+nVbR0ASMmixk92pSUPs
9eXGBv8MA7XHamfJvjLRmgA/eJUaBimUV+GrUyE81B0hyDSYT284WLvd2xioSQV3WPbnC+gKtpJR
WZ4R5516WEKIgufMxF3gYxyC2NwckmNZVav4XczG5Ixn5nTwBa+ccNrGniIYD65ACEeSNDGeoIUc
a2mGzrTg7jfeqAo8s9T+9uTNRZs7jj+Kpq1clNuU+UfuGAYWK99VjIJLB3xMtiOx6B2z4uwsOO8B
1pKKVvWkrs5ag+oruMfHjYP5+zLABiBK8u/Ve5P4Xp4TsILkrdytot40kJtEIiPh5c2bs/2mc/Cp
7zLxy1Olxn1d+Lo4YLOGRJJdtk4vHcUD/AC6kmvba464cCzciqS9SWjRaU66VC+n1b8GK+G2zJaN
tMvkfWc0abwytSf9sMyCFF4IsWhLEPxVmWAH6r7C66ze3AXqOdeTF+B1YTMAoAquTlJCjcsGZCO1
7oCzzqQRNnCBaf0hWYvLpBiXk446GhQ32dKW/cRYji4Puwid4g7ocR7+cp+bmNoBDczdh8dIOhGq
zoS1VHyZL1JdaUpqrDyvL1+fPdn3V3CEv2K2HzjpmFdQi1gbZa5Mp5KJDTKTPrrvDLq90sHF9WF+
L07CS1NR5K51q1i96P2FQQPXCTOPa5XS7jIDg68BsqTgC6AbdnLa2shAyBkqBaBpc5RK/rCVkPg/
PQV+3dB56nkBeE/TzQMySjcJNLCjIIx+3Qq/0FPu5/58xArIdb6S/7uMlFn1ixgz0IWw9sItwdMf
Vnusz6mXfqTY1C1ncBQpN/Q6QbK0P1ad3OmFhuJJtIJPOtkB1zmf69XTx25UmlTID1u7Vgt8yFIT
J4o949MWx0pUzkSB8mdK0vctYsJhkaZJGY7A1b3dAKGzuj5V1rY5J3x9ydfdgJZSI2ZToQWNUpz9
JmFAUy4YfrK6Kz0DRNrjKUmwC1SYgO9h1JHcrpb3zDLzE4atibZ6wD7qlB6wwlOlmQV3QT7kUZQl
9ZHohrJwQ9q/zEwa5VpAswREt24dKN2yRLBvSdLdI9SWwlPL+V/Eq/e8w/5DqjPa2vWjWhnjIt6A
sbuFeF/M0JT0wRFhI9Da9GhUsB5bz8THrSGzNvt+XsGbcPoFgLRUBLIaOZWq5FWTP/BN1fNoupVo
aPdogd00yG+2MICG0Dvw0UhVqwvHX8Ami2wEzAxLLJvrkMDuy1uZWKwcFk8qi3UnlipmwVoDPxSc
0x+3FLFgi+nZdFnfUflFCAApeUU8PsgTM/mqZnLlK6/MZMnR5wl3+/LlVwDXQq3tlJ4YOorwo+yW
7w7i5Sj6XwffYFjVE4oq+XTX9CNciBhtJLyEANkKfHzj5/Y0hqD5ZTjc+PO68qsw6FGaqbB1ti+f
6MTeEQfNXdO+D+S92riHKlINWckpCrqxkUfOnuXIrdRzJM6PKp6jo+uLhClF23Cj1HiEwBnAJY6K
ZPJ4vHoD0pZIVwLXIn1wovEyDa+5uz1rppewG5v9/CEgvI77liQCRZZGVvY+xHGD91fIyOjpsv85
JnK18mZjzyLi8s27h1QbJ1afgOnGx5SsFJhrgV4bq+Yoj10y8qCzgvzEBkU+wgCp4+Oi9LdOggRA
3h+lsGUlmBEB1zVYje5GfR/XR2VhUI8kPMevgEXHPuN0VEdPdQZPLVot4Sf1MuwPrCMK5JioZ78u
yS0FBJJgdlE/2EZQmEGRgy0UXFI1woZuJDCzCroxrgAL7MN+aH7M/ST7ROEU6iacbx4DXy0L5bPc
5FqgqYtvz9HeW4cz19tMtY9ZMe8C7oNzNvPlmW34AeGf4ZIYFkp+HRvTSyPTE0FRgJRpq5nW+jx4
JMo8L6TU008dmI5sQQZbVMXANvvAP7++4uDf4yqVlha02vlG5r7KV+oaWGKlRNHU0k/UAwiZZqET
yfJcMH7dJ8dyzPuEwxNiW6MEaYgvyzgFroesB0FQfjhBETgMmRWfEfXj8s6mYmWwq0G9zfriap5s
VC+O47mpU80jsz9JfZCbd22sEI+wFWfL+jwkFQAqWpxeHMEP+i4+zaqwp/viRseOr2H2BlvHS1rx
MLJblO6t0/Or+Gw7SFGrKy0W43sKDJtzrtK1y/37ev54z76sGQ4JjITdENHguR/sNmrR88r5NAYx
/XcqpXb0SizyGypgc1C8jBzVBkuxI7ljgDKxI6u1Ofxg7kuZcQYJjiHRwIIreQC8ZEBdFvX1eE88
BEzLeVa/ByzYKgGBo5dbpj4Yo96EJ1rO0iPGDFTeesxyYLxlyXsKc60qtcAVyvQl8VM7lXbxJncI
JJ0c5bJBYAMcY313XqY8esLVF3hmbwO/qIbUCbHVDXE+QqtDHGbem+6y5jzYs1ERb797azMAK+tx
+RhSH8u0k3khVxB+548spUoJvnBnaNEE3xaUFK0UkrhmwPyB2bxIv5It27YrAzmMGYigFBqQh1mW
qIDXz07zrixF4jDm/gWSRYcWUaY9gz05G9rxj0E6eAUzAyDa7ZlMaSYuIichp6aUIKRzyddBvqDI
7l7G9nl5MQJezy1LJiI84EXZf9lJT69YYaoVPoZL4hzfUldeD1fwJ775Ez7Ar4muPEUwHMtzthmM
O0qtJEcmID7Lpd3Swf8w7sFKCv87wAW5uEruHTGf8/4t1idzqKYdFxXyVzIPRHfFpIbmZWmc9vga
ZIb1EtOHQH7V4gRfZlZ6/XmbvgZbVhKrnoX0Lliu+E2KzW1kHXJgjglA1Vvc1SYXGIVc29hIwCxi
ysWITR3vBElaUdVUo/FCXn3fYbgq2WbP1GdCP26RCkFSZmjKSNxWw2nZlMsJLVCLYTJ7Z08H07dG
/NJgalXFM58/QjHFfHR2CPh/0xKlGobdQdCBuWqNYMsma/qh8fqUUiNlMGkEOpHJAjY1eL3zQp+v
pLssE/+l7Wle3czDrfCA+axQpIPwTsLtbXTjcEUZsmisMXihV1u2zWQFZ+LBDwqf6eULa4gHMmez
LZrviCc0F4bJdmlLt3nlNBc6XEaa/cAQDe7foJP0yulLCm+qjb3cI6E2LbgW4kslHpOpBZRoCVOm
sOrEj/5G9szNOOLGVzL5a+Tq3Xy1AqTMOmZBoASe8xrXq9mIVKoBI+QWEoD66pT0qD+IsuKhszKA
dx5ZSU+TxaPb8sHJT7neYmb7WIr1UhzLtXl33zg4dSaQdzBtAhvGyyEXhPQBvXKOjpJ2Z+3Zj08i
OtyENu0chnigV5WLnUkVDjMn2oFwzWOve0H6fiF3HXxOKvjwFDruHhwljxE9FCY0PyksjAOcBtZX
j+zh4K9QGbW8dQbp7T9vMv/3JABx/ME2oVvUE0mtknB1oLKTRfbq33AYrONkZSpX1Y5hmRPPtvpp
oKGl5PzlD8qYQ/YQH2HLBcUbEqpdTzuLOkA/nt6TykkBiZJ46AjdNgtqfEtSKjjyQZKsf7utol+n
jTc9JOCnnKLdFXc/ZmIDOYn05kO4bYV39vSuBBcq52FUjgbPUjLcXHgOyT7squMnzLhb9y9DFze2
xLykaKKu0pHJ4RZyDR8e+d7naE05Qzo4MZGKZYodOUE4D2Inh4G8raWuZ/M0jA0nK6rx9BCsdMRj
oOgs6tsjdYldjF0I5mk9iU1ZPTnLwWLbnZrdBaX5xH1LOlHW7Z0xlu3LDbvR24Zw3oscBG1reeCd
Fb0l4VfQv71TgfPUg95MQRd1g1cSqENbWBIpskocE2e80tS8J+FVTQfgVOnS0ctH29SvexKx77he
nHsGgq57IF/8cI+F2P6U2QRcbbzhQF+ajjJqYlCE7AShKCoHxp82bxkL9EEt7NMKwFep41ZrxIdz
MPU9GFVLaD2gjHdcqURAa2Ond1CLTJCUi9QpmsSwHzzdxN4/0Q7o2fNl55LchdsQQ+380KcDTGYN
flritzih8wyp6SceqUPxbK9ZSq7yN2HqxmHda9NsLSgY5L6Lo7yoI1RQl52ay7LidAOmU5yIgQv+
OlVissGN7SmwTcdc1Vty4cNlUGHo1pdWgHuZeLn1mGs3CQWrRqxqvCWqpi0pQ1pu9jHIaHh953LG
lKO0kWzjjtHhpO81/FlqMf3eRuXYAXttUDGL094plGktGIY83aM2VQBylPWzQ0AC4M+9LauxYNRQ
jJ348I55sv9VUCqbiIkRhMIsxR/YQttb3jJLfu//iqfRs3b47ht6zbMIYey0pNEDhHp+nYX3uTs5
gX4v55qk8rLOzH9BLWAK4vJDEAgqvokdCZKOsyaoHirtRirsATcsQA6r3vHlYo5JaMMKPt73csG6
S4lIvRkcIJ2HSeXx9TVO9tncq8e/1KXDTqzuLIkWC9dV/Vpt7zGCaShBQkeb9kxUcLK6rhHnL/NE
qua3+0Q+ydpDq0lMeNzyMjBK3V+r86pP7uA1EIITcvsUC7IwCinT2n0jEk4nrIwrGxeCQtFHcRtD
G4NQV4r1H8rUV6MqJate/l6O0nt9zUlJWYauTGXcvazw1rHYYnKQi71aO+aqglUWs05lEcPmE8xq
iViVCA3aADXyIpsCFKzHRzhG8FIfhNvhFiNc1pV1+typF3ekUQ3kP1RvuKHBZrcsjaJOROdjgUwb
c0G5iuaKK7ZPFdu+lsYEhOT0W81Ng4mMgsbFwWAqamoSwYPxs2kjqo/xXXfy+fHFJN6miXr9AsOo
CaAJDzgL497Npg2zGAIfXLfuVYytLwFi/FFusM9ZBOvlNHXa+V6tU+ptIzZfuyy1j6fZIkgB2mAr
Tsb7YCPmYNbokGKUtr+Ix0m1ILF1YOxTFnvoQFsPku7R1rHJxTOpGVhXv7rO4g0sEEpME13zHuO0
rtQqrfStxE1Lgz7fI8f8XT/czq9eI+s9zKwhiyodaHQpQQiXhRrLHbQ++GAZNTiM+kC3vsgv4vhm
hjrDwNCoijeMGHyxGypVeBxUClcA3mz1ClpNeArj1RTJ/SzNN1D1lXNNRiD2U+NBZ8mgWa3YUb6K
Om/gDm9qYuEdFkWr7CoaJ8Hr5buO57WpsKJS7Ta9K4xcjRP5obEcfjTIaMPzeZy74DGInk4YfY6N
jfPRDzGWctj5MEh/ap7IdJfUUBsY5/yds5W+PIN1Ofez22u8ddKArFSw/Wol8qlQBl7zBxFbKHZa
0R4e4MHmV3w046ffs+GNyxSTRUuHTVZITwWov4JVDzOh2mZoCTkwY9/U6wqhrfm7ZaZQ5rkLtaT5
dP+k+wVjnUJmir4slmK4AJ5hg5sTwrSeVNfpX+sOcF0jV1u5D0GvoFGfvpJR96PrZ8fKbqzK4WO5
xjNW0+ammYNY1KP3sJHcNXaY23qRxx41TDsNu5mU5BMYnpgp9gx+wO6vBF6h/pwOcKCUnjiTAfjy
CW1aPEtALzyQB1MxyI8pWeGpCXWkFYlPVnHnLGHiUVWcx7fGlGFhqoUvbGfkYharKETstj0STmU3
u221uK6DwmJ3hMuHwhT/P5looH91f1pPTkGAlLklrFxuVOSJHw2Ffrcr8JJGtLS2Y9VYkpQqLsi7
fxSaz9S3hi80f2Yt2zwHndpEnILRYzAl0wDdveB5UOWfJgLAUEoYnZ6y3W8QfbVyviUC67NlqQeH
sPHrglhl+8XB27PI5wzYWvkSDmGv0J6k16OM802DjeDO1P1IMBdsL+5ELAdgIkSApD00VEURu0+6
R/MkAoYqITz2L57zRSMVVX+AyoUBb8p6lcFQFUIZWdxSuVBfd6wUmkxT43gEN21EYOvt1kcF5Wrd
dHv4ylkqk1cYlitCYI7T5yTMIYFD+L2z9qWZKc63Z+f60Bp/lXoq/oDO6Ew9w4bQJ3Z3YcjSb66j
dC/aHkM2xYkvCdJ58H1jChE3VzEcEAonJCXJbbcYaM6S5N9R1NVg4vbicAWdGtLYj0kr/JjcAiod
VAM4zUIQdlX3sHUIp3zSSqnZxeHSrw/5GLLG7IvX+o89RcexsuA0+2011fdYnWd/k3lrOMB/OUZQ
v7CCDVLQK3P+ngRsGQndsKpouVJ92I7l27lOGAF3rcAxBSQVZvsv0SWEvz8aKlILIs8GIwTDDeHG
pxld4yhbyqHRwcnMYyBo3Nw3+7FOhnQcMhKi8z4ffNwXCRFXh0SEEDeCMM9t6bGCa+bEYjwRSMpf
1uTb0vvo0hyvl8OEFRDnCXmaxbfDQwfn8kujZq4iaohj2A+Whxcx5tT+At5Ex+L7AJJ2thIQ1cKi
KFH7llLJekKTr87uOkF29U51w7EpL+mv2tMLeWm9XaRLeP24MmbGsrGy/eRv9XtPyJuCe1qOLsk1
ljzfdovxz3l0t87SQ7wId9OOjLg20xce8kAlUvWQH0XNioVgmi9vRVMCjsMUd1iKTNQQaFGBBqOU
dilKrCJLd4y1GQbFVuNC9iD9yH2L7WBuBNJ18iphJOHbu9bcmqal83Q/9mh8vD7CqZ/W2jpPIZ+1
5rzKNSO/m2AB9S8m16asxG8MhAmYSH3XeqpllTeA3+TeQaxj8+QFLysXvWdsswleLN6GQF7wYtSe
L1h60KG2MUPYLqhtXSAZMbFYBDS11A3Br9ecztmb/8ODfX7AX4v7TwpV6OUp4yBKJ/Iae52Eo1Lw
LWJSboRnAyNBxpOmeTgTN0XYecoaLZF4Zc8w3SLLSNkIqVRCWO1d9jttOl4Ljf4EhpNK2BbKjTyB
2EAMZPHcDhT7s89+WYrl8ccXLyX6TEiO90jTkBqxaHJsJorgihVosMo7eWWvL0u4aMIIyiJgw/uu
2ljlvGzwV6pytopw+SgTBw1tcR5plO6JrJFC7lnNgu3Lj1RjKT+NJdRXIsD4o3CwhWzk0wkxAqY6
88i2WjdoHGYdhUCzcQuROVO0UlBTf+4BPz3jtk6gVR8fLGcaUnSUJWHoolTh8DgKewKhq7bf30fZ
JVgMcAhq8ulb4pECMKzFJ1JDnEKlsnF4b4iRb5wuzXveETI1NDu4TJM/08jTrafUAaT+MaWDI4Mg
9xktV91Wxo+62CH9RwxVgPnOMdeT+hc8L5KULCFsmboQOTR/bURon5rihglsPjwANVlKRgrKtWgC
c2aRl1DvW6yAf2FrrXH351MvoFZRzu1FjNJmvE4EE1IrG8Cj3c1TNhzey1gDQaJk12Cs32zTloFw
NK5uGERPU46g7Nt1i86VkDP19zPLmRHg7csd02Ii4L9KL/UbcolgA9gStWfUYWTKr4vSMI1aDuRr
RHe/CtBGT6u+3xJRjk2X1xKahv24HnWMQQs9RuDYE6HHKA2LoOpDGInXFOffNbKrSANSP+EH+9FL
GS+GtiPYv9j4PM8TBA2nHE+j2y1PpGEk7PW4TuxKaIWnNatBZoTh6UAHqIv51jA+Zb798PV5DbA0
c9Wfh9lAbawDgZQDruW8Zi4cAqpppwJTlbOdA8TsDQiAjmhFj7uTF8exICzWA+17KxW4kQj9EAAa
FpFt6ijI0JpW7OT6WCDOPkWYUbdyZQtA6L+gsg0RFt+ZmPN1fujq9YB3Rff4tr2UJXm9XnnEVUDv
SB5oPgP0Lphh0Lg8wjzqnnTmKroDr2QGQytz44D9lQeQ13DhbFiUf69qu5K05JY5Ejn747jf9IKi
d3/r3UjMg16hS4PdvLUNa6wwCk+cnRmHL0Hi6n4CB8yYb6ncyshqJ5zWSNi0O/qJSWqJ4p7Di1oM
52d4yCX2Gs5WDiIR/fiMDW+b5eDBw+iU8j3tRSHuzO6ZAmzRXUZ9ShFVBZqkr/r+1mhPVpiwAK2K
NMlTULy3ywGOtww1ysStyKmBfDpI8XDcyGl0oAuVnOjnVN2q96U7TnYJoTEWZiVP7cVb5YY5a3fF
b9QyAxAfdi2OQGmuxPF7NRr0E692zz9Qxvq9QFjYV5K93d1Wc7sfwXWaoVa/Lhp1pX9iiSq5Wh+f
+Nc9kah9Wzc2GKmrPTgMkb1HgPvAVX7Z4W3mmhCdpQZQEPbbZHeW9RDzwvtcIMzTAHPxI50VoB5V
yl061IILDPLTztK0Uexxw6+43p5Qy4LSUt3u8NYwj6is/5GL4dtd4fnn++mHDk2mz2HJ7NnhLLzY
8RRaLwDmbbrooAMIdKuZJKGrJ7fv06tTHsQ7xHvmLk44rPdV5N7dwK4suRmfTnmNMyTyjgYFf8S9
3ct2UNYUpxypJ5tAdNksmuyLxN+lCHVMyEvcGf7L+hK+BoVmvEm3RVhCMLl0/Y6t43ji8eJYOWgu
g43LSHWDN6yu+bd0N/Np7v4mbS5EKRfV+WGNKtsaGcmUdUtYVwsb664DFm2T8k7j3NYdZgsfjhjR
6zpqIBjD43ykk88mRNh7IT7nOrTCD+vtakNL6J7urq37YvTed4XdyF+9zs/v8dqYC1Bt8hrFPYvS
xDPxEc2g2+wG8CiCwWXhWKAY3i9IyV0su3j4RPyehM5t2qXksJ9G6/2OobAnXDeZyoND6F/+1xnt
0v+FPPhl6LOQadbsmd/BWiMK8ISb7jmrkGHUCQdurz6uxcoLJGFSfhx/7uGyeAa6S0z5nzw839aX
058wamtAFZ26840em3gYTQ3vaCPP7AJlDo189jzZfA7Q9RdnATjUhJOAnFNlxToUbCHE594gssnW
Exw2hJerKeGyG9r0fNERqoKL+Ir2yEYrPTs+MS33JOzVoAi2cebxMjYg4Oq0rHAwRSmOCd/IzndD
tqPyH3t1wkMNTqEMAgAR0uxU0W5LTmJRvhywSzsMZCk/L5ZGErrwCE9HR9zxyBYQUP4w/ChwfWKT
NG21Smxf5WWYugwPCcNYmHqXsILlZeFxh4nDyNipbXFvwq0CDyaZF2yYA/Xpto2lfEm4BgloUpgR
LtkzimYbP/e+EzO+Jr7qd+5mdOMHATVw9qxlle1UsC6vsYNEaf6D/1BStFZyl/RO1Wt3Rjvw5ZNE
O8YBnbLPOmpgMWtMnGdrBRKjoAGHhkrdE5xVtztvkaai6Ytxaf91B7hp1EmXEpQuWj0zyESwvOcs
7swzhFnfjjisD+vZOUpVgFzHjtFoy6mCr+zeuywUUps4e2SWlPd1ImCllq0/qIlZpV5ae0UYqJsH
FtQ2LdG5ic75eMaW6jQrAT5wwKJQsOS7ogLzBc5z26gcR8GD8o3eToNXtGQvxmGGm6AAhKa4ykxF
l0dwPGsJuOjGx3ythsrSWQRf6P3EI6MjW2oxO+vpcKGYzNMfN9xLqliuZJCifA9CpmcOazaqDa+I
gdsKvTkRC+L1lJx3MYhdX8XoEzewWOYS8RiGCd11whc33TXSbSKtYnV8laAi8fOnsrxLwid1FjeA
usag6UhHZENqws+YMujkoopA5UmWqd9Ytb+fDRn4GlNpB6Ky/GF4oM13sE2dUaM2EQwJ5tCgzLJq
EoKrY6kdse2WeohlJz7M+lHFzRmepNFAhMTBgEYWkcT20fL50UGcug7O0aAqKaLDZ9a0BadjtFd2
RVz59f5aD7XpR01+RG5H9Y/Z8v3bKdydEQGuucE+S8FNepjFGiFL15JC+15cKjlyKaqp6sX87IFA
1cD9egxbhT5fzhn3oar2r7GQ+gKFPrB9azF4aE5yCC8wz+Wsx8Zyx8uqKl9rkpjWUrcNUqDLOUxh
o6TTsRQddtdyeceO9tKV2ir/0uUgHxqSevmMu/rEIfcoLhTLXA0K1G6eDf65PMwsUzDxQUAHtWI6
Twda+CkS7TpixtotAhfB/09xxEkBE6xoPET7hXGCBbstN6p1achJ6f01jd34HjQJBvi3gQ5lZaFk
1rRN3MGoHKI0NBuraZa09vDOj6xvbD9lVcdOFspxQssiEd6Q5LY/gTqJLQYI57g+a2QvQliZrjhF
C3VNJF+Uq27Fap9xJy72LYyLajaBLjVULYM3vwtYYu0mBgCI8zSTh9JR835H/KTLG9pFfo+U5tTN
/4vwRe7DNrfuTb59RtC2COxTdI4oVQAR5+YyaXy+dRV6PR4qmcpopwx+hu00WHZYjGaHGf+Hs1up
rfX6DcmWQSwp44RacK8Ba5uyZUNgPq1+MyGS7RZjwfaRMriWfvQaYyxxxG+S08buo3duC90R8k2V
5eiMNegaFr8yXrEiWdcIgotXuUkFPrLyGi6R369mj6eaAw3gdJTJN/XJtrRWx92LNRS9TjaGzUhU
FepJj74i50kwBvdilJHae2UcUnCzm+XvaMN80d/+Bi086hMVULvjseE1+hTyB6pzIhrvNmqWusPu
tMTSVkjNbJCUchGJyIQUGBkxjCFT/XpclWlOCbbbYLLpm48oTG9fq/b2ZsmcsLaFdf/1rLpENkAG
D9fXgRRsmYc8leerqwAx3YwHjAXWTxy1PfM/BiChf9us4ztudBNU452tyBHfJR3iF5gfPWAvJR6Q
OXY84QPMBN5WOoy/BiBsM3YdsU+dBLlZa0Ikr4k00cyab0WQSikZLJBE9PVG5cBgF55zre9vy8bS
z9rrxqov7z2M5hd1VaMrQpOOIlnztOxqVQvIvVNTXe3XfIGVLUP3yHxTyQaRYBjaFe5vQefc6cem
FYHYG5voAkyT15iwJ+xW2kRIoPusUuYiQwizRVqr9cDVmYURxEZ8V+nGeTrzTRt7j3dCYF4XmYMt
bhYmYIgb4sGILxvEGX4ogIDZya6A8019bs7dMYBLtAo0OE98YWghKQmmB/6kQ6IABEZQFHRmQo63
ZnzIMQlPiA6yTEa3tIX1NLyVZIVW1aGrPARD/a8GAbGF/7ti+JzAAj19Tqope3qN++BnoK9atnPK
ILpUOwsEJmsH0wcjggXyRYopglwNwMsmgCA8Fvw0MR8noEzT6FlvkUFz7iSey/d0msdUuzAr86LO
Dp2JUYu6hexVdP+fY5GlNDKtOsR0nGl1YVm3XsfsLVhJym1bMjtKFKmvxe+zrKLa1xyxzH1e6YKI
FRgXou0arCGkTY8qmouOvKgxfr3QDlvWX4y0kg176vDqFd/r98F2xEfvTH0yiS4puqguD3pcI06J
cEPODEo1rdIYxZK6l+Elqq/MCidp93/sBH+SGFsKmE/0G39t5lhhDWHolOgqNyJZRrr+gBKE07Qc
6la2vF2b0ExuDrJRnTL+IeRiQ949reCDwO2/wzF4sGkjcqEDyd29nhZvaYEIuiioVJ2BukRsc1KV
PYvkNiDWRh58ns0i/RBCzljBpbAhfGtcldniRmygpililvjSTwM18BCLCIXR2wg/EGfHIFZWHDyy
kLp56Kuj6kiCHOAwrAFFOJ5/x5dBvh5aa18e79cDmm11X9IfdwBiMIKsSqcLT5MB5tnoQIKqkpKE
dXs0kPmJJcWX+zYJV6T8zOS1NWsynheShj5/j6dUaKdD+n/kf3Dbfg2hdbhr3FTdbqNcTBfdkHaM
1DJN9N9W9l3y10JlxGfJp5ddoof5EDA3YUXqgDgfwd4EGs2TOor+DD4fRmS54EoZQQyXu0ckJFTb
YIKaNyl/htXmVK6NRdieJgq+0U9xs4USEZ7xUQhPkgzIOa8mvAjyWORTvEMe6uGNb5wtpRUZlYZI
khGbiJqUeBkIu+frLheCfx2JPEa3liUFPvIo3n5Vc5v8/Ad21ddp22nOsfdKS33kZ6XTmac66Km3
KNIFVov+kPT/7IbY+Ap0uE3bcJQmjB9z8QDUWpWpJIb+9+dKFpqquUbdsmrKNHpSPLYByNLY88gf
CJlgQj4AEUVj3K9lPLAN9ntgytugJ60mQ0335vhSSYLncfXxLB7M1kivB44m/MgYKDTQWZnts6Uy
ztXTuC4b+NYRAXlLYa24ckMWYXgXnEWoQtq8vgo94lH6esm1+swjaP39/IeNIexfXwg/qc/H+8Pu
Uhz9y2xYLq0caQQ9B0JK6a0nyGKx+nNBv2pTLfErETYwkLL6MB7ZBHzCsV3dRnd+lnpsaWRpTv6T
f6A3SDNhf8gXZU2haDfutn7vUVgfOI/PgGF3Ag6Z8hTHlTrB7PEDR+5oJ8AGu1bqM4YJH1LqpfXt
mZLjkmycMhU4xgbQ2v7rYXHiWGnrdBDFy7kcmKxBUQ8UIoftx6v4hXjQX0USD9NQwZiGM5rmO6mb
X0XIE4wkXnAdOPHBVJ2QUa1s8o8LuXFPtbZ9yatLdRyIbTX5SYV2aSgvaEJTgqz//V/qGrSeg+H1
B99dhPcOblb9FLniAW+D/bbr43ZPXmKljBxWvyBiGYrO4lRc5zFahp975/wdCEtTFLxReYnXPF/U
0Naf7asJSMucDBxxrtiLnxWup3qxHEf63TZorL5A5gICs3x2Fza4sR77lHHP3vDbX71T8RhN5E3T
3akIJJtv28kTgU68y9a4k85iJ6m3bQF58ehAVcEOnijAfvhxoQTDr5/9uwyK+iOt/454k+dBaDDR
IaU8EXa11cIzfeRZCEu48tbvdXQ1Vdxwtx4GwBx4cQO7hkd47/bAhjsSXW9tPF0nKUxvCNEmUEh5
MTHGVowUP8fN/xeysvGIdkOFvF0BMHEgotQanuVn1kI8uJmJGggZ3CHBhJ6A5puOydLxbcT3DfOC
dFROH/2B3Pd8HkL3UFHj8G5pzTmwqww4zow4DZxfIgwC2M/Nk5HTIJbopD2uUaWHNcZuA0WyRhA1
US0SrZ7QHDtUcHNQ4pwM1AI3vYYqYHt61ku6RqnmfSZP+sJZuofvRXNXvrF/Q8vV2RAEeG41Wdaj
KMI9a5/hAugy3i2zgS3nYtr7YfCXStrXfwEuuL7Tbs6edxo9faZPiiYGs2DlYHBWdkeBe3Qnx/uV
SGhniK0W/HCx0LXScowtPnTMCfLO23gW2OB6mVlTkuhRDsO+nZTl8ik1lzqIB6waQAyhkalPZgtk
YYvi6IYlsIlfvjPGvoXJp4EXWy5Ms6SRhAme6C74SAdyODBE9j7QMtgVZ/5JKwxgx4pHkVmjqRsX
hOzsaMy6i+wNf08+3rZ7sT56ai5B2w0V1op+SdArRFc879aZjAIEzAbSHlajkcsuMTBcQbt0nrnQ
L/RsobI6C7186I5mTnXArshWfMHq9Hs9De44eDM=
`protect end_protected
