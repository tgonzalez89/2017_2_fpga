-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
P7RpAwfNG0/T33mmEZx8kT4pCiB7Vzpm1PEDaIyLO/AKC4+NCWZmyFJnINvPUC7wY029tpRXW3Up
BA0A4GFLq3N+JBYfnZ/UKQeOS6UbG+OosNxACBFGce12Ny6p3eLZvbpka0YkiV1kmAOuBBxUUg1e
3InU1EgfElL5ejKERb5jFixTp+aWAWH9iihPLkDJp3Nv0YP4kAXTF0SdFspI/7d9YkcOO7lJj/BF
xp1qgsPPd4f28p/1OHr147ngeVUhja/tMHoe9MuGqtvRC6o7u2T1wC15oLyI6y0G4J2qAQaS5b3Q
zRwfqI82o5vb8re0+aHR8UqFHfdId0jHiQ5yLA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 46032)
`protect data_block
1Ue9y2QYSR6gy+4boE52cWoMF1mSnRtw2G80QMXQrZw0DFRo0i3KbNwCKY+DcZBcwBXtPruQLa30
BlLenjMGxvA4JcF1PuAVtxXnpvWawIF1cSyzekwwcIvlrmOZ//Kz7DX8z6RIo2xhTIdAfjpUir7S
/3UpqW3NpB+b+DJSNrfZ1sphc5keAwWjfwH9whb6U1E2NR04IUE9Cl05/hm0OhKuvlJ/ZnrKMzUE
HTQDHdGvi/O3dFgEbpHp0c28kFyLSeDIy1q9QVKkOyt2+5oZ1QWRK8milqVVXq2TlfaoIEf7lUdz
XQB3+WRoAW7HqKU87eH+bOnl4ciVpS/hHE8wZbtvAE+76azeu8lBmqz7/Tvw3uBbQ/gt5CN8KR6t
W3hGxGq/4QCGyPlqV0FzozkzKWVLXDy8cpfKJLhcqB5ERc2rQl5NNfGsiXF4LU9PG5Ddzjw/vyzZ
h9+zUBj3gV5ew+yvR/16ndGKmjx4GtRjuuoHVXVg76N/791s5iDwJnzCE6zuNdsPW+XCTOL2WNdY
86BFSLVir9iysLIVht+/QMzLQjldKkhH0avAa+YujpKiPYqgpV0iywCG36ZW2DuAXmoxHju3ElFo
5+HTo+S4+oeYNvP/eVDzAD1madEFgBtm5MHsnVV0y7JW4z2oyH7U8JcL3UvsiqOyq8RVdb03F8lu
jvcVG6FEfoBSqkU+uoAu5HcDz+tc0qVsV/59Brkfc0yTpF42coDmTyL/GUcZIyZjxesS9p/eqUcj
zlEVZXueQste/ypZFZuQwNu9CKEC9AOfV6CurGxU6scpcJrvY3Hhp7AY769pSNdk4OvE8RvH6f8S
OxJUox3nOnbGT6LdFDfapsTEhF7iLBEScsJG32oECePgu7SGaq2vWPy5/0SULNHyN46Hm+x7g/Ac
ArYp6XPdLR3irIQBSsAYxuZi0CqVR6VaYwHiXtqTn8eVJLO911YxXUn0xpuDouYVYIvSkmh9p2yA
m/OLcck9I3/tUMXH3msfiv5glJHEtpaWqF0ristIs8OdJuMcDg31BiBoxJDgDlbasahFkcE6ppDx
TSDm96iRWm21p0Cj0pMnFUpWqyTwXqwUvbtNvZuzRuUMmFTyEXAjhfD9K6Hb32T3rIO1jtHq3qUk
Z633VZS6zM9IxzwmKPd7FDAfkbYgjJEBeNNjBb35LL7A2NhXCKu2fALWwE0+I7O0dnBP7kPZmsCk
UXfpdFDl3YGuY2/Vq6Zj8qqbPnuDn5nTFhhKaEM5V1ylyGbIEBWmPChzmbvUIPGoMxSMoAHLOEES
zCm7KFmUaAl2e31lzPQ93KtP/f7yKNjsjmZFgVodyDPTAZwwHFYN4VgUAy+ou2vMPOvS0k7Il+NL
YkJGX8eBax/R5HXcTpUmcrlu5Buc5pFnDPQbwyYo6einrLN1TnoOKzOGIMgVMYve5geOGBoaPC3j
fde8B9RxtZztmLqHU9w5LhlW1n1m34bXdXDvs7EOdw51OeljbW1LWv/mltEL6+Mr384q0wvwn3FT
mTTodjGUbtPsVhWObsNFO7tig2D/XKTUWaoQgNrnZBoDkFkKqRv9kcuThwsqZ2YOZCtz97g/NJzR
uQlM9kN/euuLvZbMSEFLUtQuDnNnIQqkDVcLTRhIcUA0AfAmkrd5sjCGVVqP69sZ55inMG2UaAzm
3Rm7uiI3xtu6YY+FHCpQZUa8FfMFCKkO/Q/77DNsClShLX8woJpG1q5eXOy5A8GvVh9nYBtWIRzW
xbCs3MNZGILEbTtuMiLKQ+n2k3sutKj/787Sr5MEiuaj+vn/Nuv3V8+pWqtXzsYCU515xVCtOgIh
0IkzYURPsftCrkJ2Jmv449KEFAynMCV9rsJqDVAu0/9cVkJgFc2LgatG1CJ5HUH2AFWipOhT/xkH
6fjIuv2MVq3tUZXvtWV1/mc+VYKYOOct7+prsGQpxTvgaP0GMcTjqfG1UJPtRqG8ugRCif5Sf3pF
d3rp/I40uQncjMkZqYmnvCn4H4hVgO7OPBGrtKYG/GXIIJ2IZvzW+KMm2Tn83FCpyV0dIqu2V1JZ
8eNIwCbVMSLbqfP/roZfAuBjprpW7Wsj0v1kbjHESi6XvebW2tti/xyEymjRxaJ7QHb5N5r3X4lX
7LdEZN7Y6BdikjQNWFKddaYsfLJZfsuVa2o/Kz7iRojcPfZWDuovger9snQkTLbrBb/dSxazI4Lb
V/GTIxUP6wmih6xmA7tODzOFHFQ29m2Ng8aYt5jEAKrkWwOdOj6ueY2KTJJc1BQBKuM9bo6ZO3OS
MaFmOUyekLB4BFbKB/6X/nOaB/cGNe9yh+Q8dP3zcmWwYqd7cCGzSLFRU5UPpvZvuJRQ1fQpNIcD
EuOTOY3YN/HIkjxZRovZYdLWmX0QPP6xaP4ffwRmJXu3DrjxMgzEccjWaguDwmGJWyLa6zOMxf6v
Ea1ttjdfP4ckBDwnCO1aFQ6B0o9yzP41JuQsFQdhvAqSo7c2C0VPOGMOdWiuSbmOGn9el5flFOGQ
I3wH50FFK0wctug6V2vRXbz6urZG4NoYBvp1P834tFyl1HUgwpIOqNdUtJZk6mwdqYeBBZ2i0eqh
dbZgYNITP9GSNQBbDhSjK4pFlaq2YZdJsxuZKerDDN4qKFiiwvet3DsfBbbnUjHJqBRGG6qII0Tz
BXqs5IWPBgWHLqhYdrRI9updGRmMcHAyf+YDF9fAbIMxd1eSbZfl8mkxNHbjME8wvyGSsu8xFWCF
fkgzz7l2P3KG10yYH0BxATK0rp3X58VHGqnmoqHE5oTWf/Ls2x/VyTm7hChhdWG3q2rXki0Q8JfW
2lmKo2mGesDOimUNG0mZwMIJcnGvMrweoVrPkSTBEgiZnkZ7TrVmAHHp0hnsVD3u5wW+eiC5nGr+
NMbZ15g45+DPt1rDJKtNAqh3EHmUgbBwtguKhxj8H84UWKAd4u5WKyCl0C6P/FXX0BH2Iz+KDhWi
8oNJyXBKWZ6LKMS7iJb+cTGvEzRQobFdNYJa42z2en8IaLRdYNGDLFFIKIOa6ZDAJ76QoCxj/Czv
Dw9S1pQFzizJEdd/BFARvTXYEIUcCTi7SspNJvH3XPEEWxRflehGZbBJ+idwWojcNp2Coc2+QmFS
UNkZzHKZSBzcv0clq6f2ju0uc9rL6h41bZsTO75WCVWaPQEy2VrE2CJe34zbVW80eWlYoUmgsZxK
CHMOn/Smo3EZI58c/4KyqBo45bcYIfW9Jyk1zE0PpVT2SJSwpqUjR+qDq4IJ4Niro83C24pu9wAz
PuiX086rwimtyn2pYeiMpF3yMqBhw44JX1iulUiKTAu249YGY/jNC4O6HCmPToP2NJHlfdiX4Egg
nytM6Mg5F+UUI1hjqGefy99e1HU3ELFA19GSLjRYrPfBKDqe54Cch6lbaTyG/lDG+vL/ewzBMCxR
PSvpmXExypb1Hl0GJq3yiWPjqZ3gKfNcToRJTMvPMO+wdxaod9oR5nY48VQlPIiOw76kSFpaChor
1dRBCb0/tWlGO6RsYJUAhgMRSfioVo+OZGPvI+hj/msV3y865tFxIrxZxbpaYSqSN0KCwnqG7Oyx
F50innT/NsVK3KaumejZojdjYmuPW2vwdgT9Qp1VCxSUSUM1sAe9PbecKDqx1csx7ep7cai7dmYV
8yfGFYEFY5FGGlnX0fouAQ6HhzaPT4y5Rwpdv/rz0DjxSnGlS/Aga0K6D7VYYZ4pc8kq3wMSYQWZ
+WNwAjsLK5iZlwII41Pf3YgeCumAQIsXZh/NNPPusGF/wHk3VDZbRRhavlbPHv4gQH2YoWKvc6Ya
pG0tPs+UNlXD8Etc3FpNcFnLxr0PuuSQkaCToCctbDmp5vzOn87KGra6E2zfFa2U7S1Kzrhg7t2r
xfN1e/fA5na9CU+9ZsKhO9fgha2t8hus5euzNu3/+pI+miX+MJHoQKOM7dPkteGX8YhvFUHR2fLr
yFQLYzPqh/165PTe+SqXIEJE7EXoqrG3vsMPCsDK94DweknXsYNCLoiPm4KiUKEQdm8/MppeogBI
E5UcmERH6CCSuzBZXr5qNXrchN6eadZ3IHrzlXKCy/Y+7H1mKL0FtzsT4pao1rhNqmUXdKLphnyT
H04F1cWY5UqCxp+tUaAt2pR4EPMS2JAwEramEDtRSkpF4PG6acc68MHfzuVvkzqSt+BRnlHOsekq
ysucsSLorseHADs8WcECssP2/OHD1NmgKhfd/AyjhnFbegYsZW32OFd3E+IkVEk3j+VXmlb8L0UW
I7k4e50QPrJlwaFjAppRfP8oxLljuuYT8dhqf7zAgGKmqtCDdKZfZz9lSxtpZoi+I23djVHaTkGz
ju/QTURaGcV6JM0xl00y/kEZjezWfgUxc5oQV6KArJuiPjavg2jfZ0s+J3pmu3JGjWW+vj4wQH9q
U4TDuv3asF0GUKZBlv6zlZ+/ruJnJrdWAhsGoAk02+EyOYsTtG9IykC4cyywAc80a4IGVJslCREx
QmUpbyS0xEuesPuBvTRU0sk1PZrl2EcjvX7Dfq4WpkFalvi1+p9ZKHdECkLG3Kg40Bu+9Fvmp6wk
676KQeZzl/41j0cUCX71KW3X/W6VoCCf6GGeozVtzNGfybAEz9fK1wFDWUaPICZdGW+ckRRrBiN5
i3L1lFfo6z+5QYACjlOATwP01l4wjmmPCBspVfS89kZNNYwryObtcWYzysE84zHXwog3MtpaWWcx
IQfReOycWzCXwWQhHLnvE7ySqreTce78/MYCGd50FY0i3hevXJF6na1/Rn6wjAqbV93SVDFHMJy+
PcM/fu48DjiK2lrUIWXkIKCTjNXuQtoT2lAlKk1YmGhGNjs1b68JX3/knBCKPP1nsq13nX+Waw+s
eH++N4eYzv8h20JiqpEakDfrh7YDTwxd2iTns7MFfGL0yth60296HKaWtYZIwqFUpjMZoAP7VMum
AyMsyg7v9JFJJBrrgAK1x/Ui88pBxP0EbtDpxR9JI9jTkdRDk1Qpr6aBiEJq/VwLYLRtZDB905aG
vt+Hqdur88fhoiw57ZTm6Bq1+4yxKAkiew4Eogar5ff/hawNj3+4G2GtaqKN/x82SkOF7AkyfFyz
q8tfEeFiWGlepPOijHd+FEEW41KYY3HZvox1hXzCuz+rjW6iDP5cs4SM7Yrsb3RdUJrOqX1pC+Ac
Ki7ExR+lw8c/yryxJA8g3MB+zYR53eluxs/i0XFI7z1oCkRKSKZDEMiRjharG4FyUZZUOy1KelsN
MY5SH6D5z6DU6V4CUvLXHb2X3h40yilEm3wXpoeZFO7pZPNb3RgwRZbw4K8X6O0GGDSe15l7Z4aa
y2ItnF0XHyKwpwQnzfiECdlH6W+h3tj1gQtkUGjrI4vZRo1KzGIF2n/RdaLg2h15bVCm7oF6Z03Z
rWMj8h7ovC9pLKqdfRuyq47m9pVwRCNKP3xKKhuQ0lBsMK+X8pIO8o/cNTpjAJxHDrB3f1XNtX49
85iadubWIRwrt9vv7acHwXcP6i5t3Is2n5G1SGP4/lJK3vTH5a9IewdRz7h9A31oWI9xfKRRWyzV
JNMWJ8YYBHmtpZsBKriXwk4fuWw8uoHx6gSUIyagPO/YDfPYUoBVPM6vqntRdDx9xdWGugU0NMgE
1Z9uETJCLMScnT7TfSlxsiamiO5TjadNV/UkdC30T8pSGvfQ5bL8nHrbc5WeADNsq1IFl6Gm+pc7
ovRNXQCAwazX7dhB0NjXH1cUtR6MAOJt5m5WIyAQ9/5fnz4k2+XJSHII/uM6JFYc6nTpgDx78IFP
gN/1oTLwIoSCZu19wLkzds2E7kQ8njD1zb4nn5ZBuP1N+TFHJL5lCJDBHumuiPNfLL4pXYtHOcfG
qALUm9mGcB1IHBllowt5wqD4eZCiO94yuDaGfAL7FaVshO7gdqjxDqLUIyxr+coGMK5FNZoSSgi1
47W7+3dN+a3/p9b4u7jX97cISyxlIFx+cVQsZ953CLiBkiSYiTneTb7qR2xK6RBd54BA+EnEFkqP
IUEiaXvAfqYmrqxsPcpJYKX8mF7Xi1w3XO4yHpkKNM8qh+zRp7Sj6kWDBzvzFAbhw3insNa2HAgC
KKjTIBreWtYzJlSVy2TtP7TXvBNh/V4Aw0nbZw693ionLigS2zpV4DUWfYA1AmiA5aoYY1zelf2u
x716LPXoxBjyIRQiqaO/9wsJyNR1hBWgH15Zc9bmOtxZQlUVZ76mCoonZdeq/qtdsRVlNEkO+831
19vLDe1cgSmECfaV2b036EPZUqXIHz8CN+UbR9wEDRAk4RvfQSgnYxd2+OimLZBBeAhrtDJVjjbQ
p1clMSDhxH9O0t+oFWeoBdKwCHrK2znUnFNL8YFvTL0vsrB+/HE9d7Uyo3PkzURPSoUs3NkEEuzs
ixsvODibKpla2I3NIZzNYQaa/lqEVbz5ahjiQB7PcNW1zmsDObpFVTrFhHLu92zuZjrZ/C+FdmEg
k7NNnIT2y2lMX+6xVc2i29LwbW/7WHshkCGx8MioggF5Elux3fPxkqHd/Jy9Mg/r0q+X2y5sqCBU
7eJWljjyFPKqdCBwS/8dZ1hSL4E3MRNh8YUarxq8w9FJrHAl8G8g00XXeFun+ol97XiE+fHm6soj
8BSdribt33UlIo0f15oA/cha1lV6PeXI6noRnjBMvcITeZyne5RvSkszTpn472J72NqJAfm80OxG
vXIP2oDJldzPo0zmGHxwZb8xprBDxfajfUOaalY4w1+g+C9N0uIlDp83H6DQteHHqURxZCdXeHrc
veZN1xEn+SPhZLhrUg0eBRfj6GULpZGCmadyvdT/Cff6rvVsCgB0hWBfGXQ7O/OcPHs66sklJh9o
8FW9GaH+MN3N+0vk/2rbc3e3nFD2+qe6eoZ6EcAvTZ+97cGJ7L/Z/T2SIPnNeORrVLFZWYDnDbeF
1vc1JmBvhkyBTk5wrABvIrMGgVJMm567+x63Y01AMrvFowEVXPe2LtSvxfzvMJXPQB4Spr+bCIxA
NR4AH7fJKytfI+3u/qu7YW0A+Y8M/lTohvqmrRxtCPgSmQtUnA6LDuo3YXUgXsYO+YeynJI/arSZ
14eHJztbacpiNNOGYk4kRy12whkql5M20a8rV2V0b/4jWo+Sbw2pv6TIcoT4nHJW+7YqrvUwhto4
oPg4WRdNsCeXUFFRd/+eTKUw9oIarglVF8JNQffpR8iZ+qw9ygy6cSseojFHuepEpBPsZESVl5bm
Poh8/Ljq5zMzxVvlKV9tC1z0SGt4F893QE1NosekzayPud3ZX4MEzoYbhArpd3BZynlYuTtVrcp0
P7PQdDMXDEDQZp8DOwxkGnXRsNiYAc2HYc6OqhyMRL4TzzKU+WmmqJKVyqujOlyc4IADzss2SGxD
r1KN/rh8Tih8ooE5aaVGxLTsdkQ2lZYeMZfn2KqL2xkrsAOoZ/1AYfZl6ZTDqxuf0T+blYez1tQo
I2rk+OK5J9tKCTaWapKB8eYoWVezTmmlT9Q2xuvBaPNG8iu7DaBut7/SIBKsJCw/7xcfJS+TBslN
4Ap+/xa68XxY0s1QpBmQA7Qr9RX9q8FOpshpxnhaAp7G9i6Ei5D4b0Q1T+/oiOojfHy/eBg87LFj
MuVr12yg82NfmkihwUTvaVeKdGMy9WOBUFkp5kLwzaBC81hjwKOfEmHcgyaFqBQmJg58T1c786zt
+Q288mSS0WKUEBx9Mndj6xfnz1Pj4t40CH4bqHSdvUHJfLYn7vHWhrbowpa7kgGKSAFhSKdOonxG
b784wrRnTgD3KcMVMJGM0CZY0matUXKEp9A3QvAv7N/LxO25sHZiksLVpq1N1bSiCgyXH9CdgdiD
IQ+uvcSlfXf7YVz50kwlmTM82BRiluOQFZY/JnKVHZ3AldDTuk+vbJvMum2sqgqDerU5t5M0busW
6ckwc2cWZ+pem0dw08EfgNwwAJXF47UNyUyB1vf9ysUYMVqmWZz6FCr+I+HSsOfyIxu6zcd8G52V
OCCLdiBz+Vd2T9WMeS/LO2i6qv86rn3YdcDFIoyRR4keuBVy++px2YM8VOQJPQALzBrIftv90RRj
uxtxYuJaPDpoOZZpRVHcslUBhtLZ2mQzY7etIzu4KbnbDKgJnpVN+PMEwWaH+bK3ghL1AShkioln
YshT0M/7pq5BjwXE2onZmOV8Q4KspZZ8wK78Pa1szmi4j1+3SJnoliiIIbnH0pLeotl8C0iKBXv3
9E4siZ3Hr/v2CAK7eNhfBkc1uu45JxdqUG4/sCY79dcE5Q6+CnZPBiP6stN0Aw401WdocZa7TOml
45LY93qaHuGlW9jeFuHGQaTMQJnOGtN6mjQcYOgl9jOqIw2BQKgUB/V8X7zQ1M+mBuMJA+HJPUX2
iXMkoV3PqAoAr+eKdU5mF+dZkiEVBoPY1N5Do5KYJMmOI6ybSZXKP9EjjlyUS+DGSTzEruRMhws4
KMKOY8mw/DoO7jagvsm3OVkL0TWrtaTecn8xm20sLecCv4Nj7oxKvx30K4nWLl7ZIISO9N7imRrF
eaegSNDUjZHtMsUQEqTYf6upymniF5cfHxnEBcVJOXJ/1R3bHfmVeo6jEbGYrRMFFTELd+Df2ieE
kE8SgV89IWxfrPK6AfU6+n7RpXKbszmilmSxlvttwrZRr8JR7YnYLIfUxvHql0rp4U+D/vSmRk+y
dE5x6HNWH/4uwdk9DZuinVjQ9ZtaqoUWndNZNjPcoIuvZAMWdvBf1e9ZttST3Ezraf2l5vs6REi8
CkUeeRjC5OtEQ1tcEfXmejjHq5AwtmZGHwz/HnfC7w0QdNHt174lPcXqaX/HrP9SzT6N5GXl69rY
3uyGWUUaRnm19tkaY90m663CSEsuQ4GFESFFanJ8dNsRgcdoPp908jezqVe0tFxVlocE0KIi34RF
6PU5exc/+ZtJTt9C8+A1ISjicsR0C4FKZC9l4/PNiPY3bdIm706UF7ubNLgN62COSEzoZCLgsWXR
aO1dEmdkyf9PISSBgN3P4acxYnrQVmoUwHGVIkXJLBDB/8MjZpXPBU7/cXrTkYX3y749xmfzRmGh
mRk2o3+inD9P3mgRHOWlZthn29KxNLKTTFcrDEw1fuZy9m1IUbobhc3ZtDZA4RV7UbyxIFR9wRrh
yx6LtXWwGhUQ6gb789jOZlKaMp/YuNPIeblI0Aw4aG4BEeWZXg/9S1PidpKo76SMoe6oohC5B/tW
InE3Al4tvUNQzh1zfZ5W7uALmCcG5WAwHEShhTghmOPntqVrREyLddewS9GmjWlUXLFR8TfHnOBo
EVRhIPpcnjcVNSLvy5SZrWeo7RdBCSu6plKWwS8Wc0756y3bvZg67rPAcAyoqBR9obCnF1ucjNfQ
Aerz2ANgn7pbOBq99vNwuqMSmSdyNEZx0qHaCpBamuiRAFIDtSdtSYryBbGiTmTY6CtrPQgG7w6V
cnHraGfhyAIAIkcVtiaHKd3ee9jCS3iQGAZHs/uP1huKT0YwWoM6w+JifDSDRiPMORvuwRD5qs4r
Mkn7FnPS2/nugBrDtpPo7pPoyAXDlVWS7VdUXAO6Y89YscCyhySppfKaI0bp68z1QnDpAX943S5X
0Pz9q2AxIRudlQ5lOyZL3FENr2Ef0Ll8+trmr/qHcWYmqWMh6biHuVeiIBiq6DjJuWn2GcoyFs6O
YGL7u3ibLVslq7ZRIQN0VBJfmpN5Cqg5CWR5yCIgDml6iIxEsQ/ZQV1D+l4Bc/N4aDUsGKekvgUV
J+c5u1t01peaTo/LRHHo3pFH8vmPol+4uEXs/9LPf0+w1h9sV3gHfrA7XZYbeDV+3EwSNUTPtKcv
Shh4VwZHK573+znBhWC4DbwvBn8hzZQpyXzdfk/jtB93cX9x2b2kVvV+FuGzNjuppsyqiiRK+peO
9NdWi//WOdmfqBhHf/bhEkbcgoHSA2dUTPNi1BcKHxtMgwPnd5WVc+dH5M74vGMCOnkQy7f7uxCb
DdDbrxTm0I+EIwuZbMzwhM0HX00o6tQKa2AHcmqHyKMQVJ78pWjBy6DIFEmXYQ7vcwOgM6Y2TaY/
dsCeden7NTlvZaiNFs/LzPbRjgbrWOk8GLgKo2AccHM6E61+lSbfp4eX4WpiaOXzn8SPYbQ2waDP
wopY9NE1BfpcCoy5mWiqOtRcBaJQGC4Iju3sPb7VP3BmPH3jT+fNo7WYn7brcm2IqKraAkJJyG2A
9NkDZXYbOBhEvTa8woReKGfM1nKZHN/e10lWibU4zck0p59cMdn1tHAEvCZ9u/Zh//Qq3bMF8xFn
pfwWuReG/OKB4OW84uujI5uXiJXtbAW3pGwrGziSR62s2rjiDnHLLX18t5UMAf/TL2IK25wbthDn
rf4VQE4AIZXQb7ua/lr772bnEeLUD54JhMLA2ILSx1yeaQODwFWmn0+5vVHvDv/8me8WRyGan3cn
5QSB3cY3t+l/zXSILbE7tHlLDbLBNUTxp35ZCHGG/JtntvFgjPPjnccV8b4u1zxu2egZg+b7CaHJ
URc48N6iEj+/br/UUgJjYcYfBnX7Ihfk0EpTe1sPC1bYoEzxJKZY+pLJnTCPXFA1jtQNlIEDSBVh
n3BUlnqCHWZbfqBrZ8VLofqE8HQYR2r/ixsST2pTNhdeX/VSK3p9Tv31pXRjejHkMP0IbDw8EL/h
l/J2DkhGsnimeQBd8RFvmEzuvBasG4ZVNTvGOmpGosfEgnoCjyzcXu99jDx+sevmDzPyalfrclan
aYJ5xZsPK7UpBEM6GVnMIJqap6jdeNIEeZe9Yghi7a2Lg+A/c1hdayerVM7F8k46wZAqFiJ16sWQ
kH1gWbWXuXYTvgBJYukETogt7obsFRVljS0WHrrSfWZsl0uUdvqjIJoreWxbTJodsVVh06wHT1II
kB6sdJ88uQGbiHK7B0aycRaONRoPPxdD+AJ5bRq180jVoDID5a4LkuoBv1xxBR4PR1gHy6k01d8B
M48tKeKnOzawf1sOOuOAOF5A2PQGDUP/DRB64o4w16VXKd3IzZBnUQAMZ6zvRt5dJ5kmZCGBGMyz
NO58c0R5sgzQIsGHm4AhOyDB08+5lNhlFYZM1vqzHLfurcYqo/C90leq7ShDbP2irgnfNKLEfMy7
3M/ZptydemFJzzc9lJkO5c0IP2sINpJEbZJcmuO1ormYa1OTTu6eL3zHPfOEIi2wRBJKiEM+Uyy/
In6CUUarMwqdLeXysjSYEwJWkFY7yL8HCPITdfvr9rUhhxD+pPlH5STvto6BpcRbPH0aaryzqWA5
HDWVxnd/++XgXfJ4SCuEaJVRUx8e15rvYj6lyZawPVopTHNZMlXxlAfW+xd2WL8/jvNR6R+FdiPA
vMD3m1umaUnzh73S3KhGgBmyaj6SkyhQsbD5fsO4yI8LMwyxgnQdxkuShw4LxK3qu1LT4MMs8IHx
+hjAw6Z6QOV/nst4NR4KlfPpQKO6qhyhjxmDX4vapVWfCygrgx+LWEkWUCa24BpLxtxx9HdJ5aVD
aaF4qEZNvSQmREM47JD9FaW1ZTgAlQD5dSXDHVcxyaoqbkOCD3HOFZBScuAIaMBSvVttoqUMK2zs
bEN7gbD59Jq13pnTRqHsKxR8vaEuzwyuJ3hvooru82QOrRh90+XMe4sTGrjCMQQiz4rCbU4nIsmr
wuO/HGWvIPYZ5jTwQYgVCJIFLE7HD8qnL92sOhpvePt6iYa7ri3Axy+NkLU/NMGL/Vqpz74eZRSY
TjVMhRdBzDjgjb74UKAd+vWIkGM7z8cy1ai7qnOEmU0Ekv8o/3U6TNepBGfQ4uxXYC9YvB1vI82G
kUtjnQknbQwy++5/p0xQ62wOhvpLh+bcisPuSlUKUlla5r7IpTJdVcPnzs/290Xkn2jUX7UdSTap
rSBXjJmfB260NhRpdpAi5QN8LIhDwzy0kYGeRGHFWH5oAHYJFqUAUe4JWTKj352YSWSgPGdev3qJ
xbcPh9BnoAtNGmMb50VMi7+wGeInKLjjMAPwikPAjfDcMYsaHRQLVTAGAn97SSCv1WeipBqJYj+j
e0no1KoULrbvLVAZrIK6/x3TlYUs3Fv4E78hKS8tM0s+vR0Fi+1V6VrpYl4TqqGgMaLaNtd5D9zG
i0ChDGH0sJtKIBTIx+L/lBDG3sM5GYvX5ddLpTsxhhF1t5vU9SQ2VGH5/Arf6Uel5YKtyEXUA9Th
G5zIdUbKUmAW2vwDdNWQSvHVyQH5G3kI4uQW4i5jYAruHIwQkkVvdIJPge7+ct9Z+xH50naYTl9M
gff6v0xHCwcK+AEGB3xROh7483JZQSizFCNqQeVbZWEA2Y3bax9eYv4xLy+0RawARh64fU3QCHYq
8vpgGAQU45LkBfl/1Iyrl40w4D/yBfj6IpHJwexc1lf4Fq23T73Ua+3vPvmbSUVU0ZN0ol915ZIt
JBBN9wStEyTNxeBKPsTKoJoZYiyhnR7KK3aWi/ntdIfgUI/zy8Yl8vqYLSbBWC5UB2PjUQhfxeZp
x1h96lPpZMyiQO2yOp6SEVN6m/P0lkiVwgwM6nmLPXoRd68pw+jkh3FCJgm34qUQh18xThgTjMQs
yuEkv0uO7L1WfqMJzhiJIvaml8zk5U+HBEQ0au1zKv/lidH4KSPI7Fj1H42YKUuxqnrRDut/VQEd
1twKnCe+f1MUGoMCJ+V5pb+xQhWk7rv6fqKoGTnozYQtJ/YxOQHKymbaexhQMEKqV+7X/n/hXJhR
geOjIm2g+qsu+ralBeH1fCckDJzTxujjV0lCsus477qQ4VYFHiVqMTHQHrCQLCfSxqpETpcGv4GI
MehlnMTJcu8264wkTHwHxKEgkyuX3lIsqq8ava2QlHirpjZr+LQlsqiCNSb695UdR6crk2Torjcn
a7jtmbpYnSaHq0L5bd1DQu74bkgHQ3uCf/gHB/NoVw5N8LhDP6oQ6vH6wBtw1kckmDdxSAZnQaVJ
EwlqXNXwOxwBt1IgIsm3GqgMplgiQq12N67PBixzky4UgnhTAmwlvCBudsF1oZbixNGGfriD9mXx
l1oZWN4uxiWB55/st/Z6uJipEE0omHdaeOzrwmUzZSMXqQ1L9EjenIgBjrLX+ZFp4gGXCOHvBd4j
DTm4pRFCKTYH5yCvCIo0XetYW2hpgFE0UJGYgUQ5u9U/Z1UHN2RBz0SIRuLjsK1y5730/v9DzTLH
8ZHuHrRx/sLxP6m8k96EcrcfTFkcCzA+WhqBBx65PLBFXObTC1YP3vWbiDsBCTXHEG5R3DxIXTUY
SjcHgmgAZLtTcyw7PyGqnyTYN4rkWYydyMvv9AoqAUZSCtAcIQD8Lcl2N+z9UjIbf7kVRUQ5A4P8
hOzzjNzMbS3UhW/aAkaVY6lvDlwWScvgtZg2nYkij02g4KAtt7bT89ny8fUGoOEYiinTz+PLMqCR
Ws9un58BtQ8T/zpWGQkUKqY4bHNqxwNSKYSrUWoPTig2ZDt7AbO6wN2YkeqGs8As1pe4Nxzx1oiR
SLUe0/eHMw50vCO0PGFguny8+pC0CSRaLvZBQq5/lr0m1inW57x3z8K1e7ePDOd7eU9IJ5obGnG0
nf/y29lvZPrModVOwVZm7JOt2AI88CJ5MH6GZLP/P27jQKUhFdVmhpHX2lTzCy/Vk0tHB9a3TKdw
kQi0l1admJ6Sp5ivhR26fBV6641/xTHQIYviXDpAsbGWa4jpA7ynIz6LD3rzE69Qyl19uuT//Nd6
Tiw5tkZfNavYu7gg7zFcexawmv+UNUSibOzWHAtDRTcPH25TEPXb1IAlEWO2hJ1xpZn/w4ydnbjo
XPq/Y/UQwDcwNUFtPz2AgfEOkex9itYVzujJC3mnq0ajT7jEauLEomAHiVj1pRQuaYTUEZ0opl1P
UZar8eIrqkiPS8X00W20VTh8xaHAo5NUoalgev5B+wrE8CwUukCXrnVCqaHfR9NypboWm5sy0IQA
cKEgwtlwGvQp120v4yNxlWJ1zq78LWLB3ROspfzHhoyrH0U9RbLklCVz3BYEdiGs/GC8bjW7PH7z
vZXKdS7SMdx49yXo9PFa4JJIaJT3d0zSVmBmRrQkR1vWlaGv0199ezCvvHH3dtbIVQgLP6Hk+C3m
8+AdRVOR7JQ0PpqvQ3XW821FqqEeprPEbmWG804zuxou94RZ7xWPErUL4LLZkXPgfI65jRv+O3KJ
5x17PCWYpWAHQQdVuW1YaQlErZKLYOmswwW2+uxJ9lk+UFeqtzq2p5oMQoGxQz9zSLo2wblSGgRG
Ryean4MGUpfVtaCSnCEE4gVLyyMRdNpiVQBlTG+VNOhac4Bpq1QIXtn9VBiMJM+0cAr5qRmakQ47
FvUAMd1a5Mds6zXxrYeTRog777YiXkRIFk5UWW2NerS99JiJ1fDbullDy1iAVqo3ZSt7h5nxpmkY
v19B3CgCx3nyGpVXNcF3gLmMrXZYsmQueIhu8MOLijGruS7+3xv47j9jO9fkUc4+g0EiKRU0jcXO
3BE4sowUWgCmxypmZmIGfjtWkuPqhQUEIhy1zaxRFKaCLqIXtKNGcltqJv2z9ln4eZOI1P5EpA1h
leHyj8a1SUrrYxdASGAsNFf4T7MoND65aVsQNWpzV9eCPT+3HrfdP9ZgcuftpjodOYYNkc3UFa3c
fBoQLBBgDYVrPde7JGxBwxll8dh/mpUIGXdRT/RaTjlGKsy5kFZbVT6oN/56cvnB1Ml7m54UkDjA
we+HNUZKb0GmtMc4Ia6LX/vaK6rBY2TZv2B8r5OhRdprKkQ7716npHJbCJHfMfy55kyzjnnhw3AP
VjKVSpIcuwQ8PhJOfLYt0g6moZnS61qbxT7HmaA6m9g3tzDQLaxC6gJY/OEEzAPUtJrE5Aw9Oom0
bD/XO7Sl2BULk4czCbtd07255XQJNZf9DtjF02c9OUToBl6sbFweV8wTMTmmZLtE91pifWLXpBPt
H5mzSzaKmuQ3c44i5Viqm7EhzurkCvZzUA23da/psgMOc99He1UBRi6OY2WWcfcVelao+eSMGenJ
z4j0kI9YmzUbI+V0BVswQx5UMjGoGmIOBgE4zNMcqvtBPaPmMpl0PW5nSOxAiKPyx6tLwKMl23or
1p6w+u56G7Hkq8ydBM4fmMmZBwrVfwWRxd7pKFnfDMuMab6MTuzoyu/HJn92/ev3T1mnkk9UKK3H
tQBoZcXV9DwgeB8bHUIjY4ykvaMSbvAOhoICKpJ0Whjs57zNqBd4O4J5dUb4z+HKd7sktaPCh7pa
S0OO4YP6Ra0Pl6LGPI/H5jjCXWGP9xr1Fukoqpc71eGNlq16Y/k6Cmm5P0y9n+EgZvTovqV0DyyG
3RYUqiNTMt8+cj+qYAoWvmqJ28p1KHxZUxSW7X+1VcihP7A6DP2DLso+99IldUWwQN0/AF10Y3Ei
BN/i650QMvWaucQLyTMr9/ZOqnyl0BxtiydqR304WuFKJQlcInRg4ZAyFDM9va/ovJOFcRD73Tge
I04vl2Eg9GIFXD4FQZ07QBk1N87haBX/KeJI6VLsXccntpIZTIaQ8wO0mvr7YCijyacy9d9ltuA/
59iS20Bu1o/BAWbp+BeoelBYpo5vfyusj7K1xjkRqDi2I/WuGbI+MvIb3xiBiOp5E3tFdnAM8Mq2
MZ9chI3YVy1BVTGASnOpNIOhrDMhrirMF6lWVm4ZHWwNJ0a/c6mv02JstqzW62wQo2QOmGg5sLSb
3WyrFClsDoX1+OVM7S3oPLQ15Pn3i58cY0MzMfKrWfUy8psSbm0ywd5mXCq3KtIpXryP3S0+ivnE
C4cJSeznBnhRRvy9Q764Sb4IKoNGH355ShA+k2RANTz+gLeYxGXyzgGka7LNGFftwM0Jd8Dza45P
m9capLUDIGSamMxHCHyDnX6ngXc9FgP2zGPif+6Cv9+Wj68K/zoawMEHw0NvzPycXZvExCYaa4Wj
2TP9M0XWMJkI6jbzKmRmyMr1dZ3HzeQLfWYz8PHSpQ/1cd7OeLsLntopCnV6ZW9UsTClShhqnGM9
zvzKHfqLSM658/DQ0J5HEWSivWaCxMPgrkAXOiyC8gOOTJjn1I8ALQBEIH8O8Sl7GOLwo7BCr2GL
/qz9FztFIdOBdm9BchKZClJzrGO+cPBfC0nUhMMTCIJ+aoxtCZu0QLp0DJxHoP15WmKLgrQhmS3t
r+am/gAe+vinkmcjcHTPAT0pcZbHwoCelzgOSEm3qVoNc2Mp04YGxY55AaB5XObBrvAADyyS3YSy
rJjIayvRg4CQpDgRKU//69+2K4/BSI2g9PY51n+yYy3N3888JlPbAcdty5+RlRBSgBw2td/i7dk0
zZBI0rVzsOldQiZbhY67+kS/XeU7NcRP5sibWoZjZ/vTMEeEfapXP3OApN6xD6QjbgL76KFDal75
cGlFXzo9tR5GtRigYxKbZYqOF+7pEyHqD9lGzzJsakiRWgCJR1VoI4hYWva4RAklkhfWfW6NAslw
bCgZdZKMn9H5Kd+Is2T+bQdsPzZXysbJGoYgwcXquedel6/+Z8M9t836aVImP3Kh2+qkk02lz2V0
k//5CijPApeoMyf5F6msDFfaVaie2bl+0/6rdYsJXzwL0Zkegg+SqaYLKfw5lvpmjmI0AIj3Ub6g
DFfqVX+7gmiYB9viEBDSEbfjgEZJb4WVNYJq0NB79bSIbcXuvNhp7OKMxX5DPr8p2+9MxyDsujsS
KVmpG6IkqLdkNWL7IveLaX6RKD5hZxZuEXP88E+PhlAKF232PU9yE0sX/8kUE+fHlZ0fN0A0RqfI
4fIZRTWOAVa7yUukZu14TqFQ0GAK7j5VSDFDmpF6Ud/l74o1K/tWZBlEHIU8zZHYT22KA7RdcoFw
qJOMW6t/XGY+lOVP49GRiIwCYaaF8qmsYlPv3VLoPiEZIG35WTp5oQoQSB3h1vMoESmGtzjXuaAt
j/TLsKoySPxN566ULgmu6Lm/XDR1yKLgqwLUfrXqpmTND5CyKClDcdhLUUtWxleXGAPN6CNMEv1L
tdLEvXM5/4k+ajYU9zBiswmOYG6fExFPbHbKkIQ6kb32kji4B7KAEXAM8h6HDfBFBsCaoaUBhqIs
qW4mZVUj0YXsGNXSRegawna3ue9cPiyTUxLuO0sCXvCuUGntdkSsAdu9FezUQckUJPNfT3x4Db1Z
TDl9skP0TfognWQmX4cHuYYwwJKc/ZXxopRJXZ0plMLKlrlE3vcNUkEjPqvUdXffOSWai06oIktH
oAUHnSDShzp1OB1JzS8OcDQIedjXo2d2GGLfbwDc3Y3prrSafIT1yaEPoh0xzhrMjVD8kzoBN9k4
GotXdb/8v93MCnVwPDOrEHaN6S3hFUSFDCsVIc6Y0GyoaFL1TZFiFmULMclbgXSFix+P55iK5py/
KrSc+gG/UhV0ASwYEcazuc+qGWkYD5HQ8qXZy2dMBKNHXNU+g8VcbbH0LXzEnjfWviKl8PhWY8Kw
+eL/m9/Cc/sgY2coB4yMbi0LJpSyUhxSHSZPgvdobAEUpHSUY9wVat+pAGdTIuwZ18LP7kvinuOv
FeoaNhskuY73MvNzIs9RK1d/sBt2upaC5SiVno5wQG3ZBezojPmkIPZ/oxzV7/ZuuYFBip2fP1I4
R6rxbn3yuYaR9y+Az7Ds9yDh7bZDweiqbmqodq++4guXlny1JDt6iXhEFd3kM296P/XNmJETGpAZ
7iZ4Ep2SAiXSeoE3ijOnR0Guk+9r3h2KFP1uXaOj7UOvjBBC0YNzo0d253I4mImNabeYESBXzl3V
rjNOLpslvqvdEaWjugI4TOAlipS1w/V79uSzor4lFOFSZ36KQQe8GdaQsXq+9OEg48gVWv10/7mV
2ADofzum1SlRb0utRqr/sq3zrCNUh5azLpMOxWqFs4GVW9lpkPnjj7Jbox5yNcY0eMOCbOTKY/3+
GDgBCBYl0KirvOdfUO4SuTJC8GiH/xgiEcMPwtxxLMwaK+lRCD8UXPem87ddXxYrwxo1ai3gj5Vh
9GEf/zG58UVc+amlJXgQBzSQMurJLmy5DAfZRFx8j8GSooJGrP0TQF5KqJTD+NHRbDnMhg/pXTaT
HiHP5KqIJZ61h6uzCmI7rs0mGj3FzC1Pa33b8PNDTfk0rf6XyTyOx7PGhH4tiA1XhrfeZMjf9GQF
s12qVScE6A++lrVXA5wXSGZugCdvAp+jklOeeAWWsG32b8M8UuUJ+86EwkwanbS679gOAalQCj8/
EZOPQJP4mz6ohHQ7RQoLIrutBf6EL/UELLusiiRlemlEyrw10tIPquV2Bxi/j+B3rkEOPIxc0Bsp
eDwQfHzBDzhoYAx2u/AelYUi/qTmrHUNbru6d3MY9jfXtzMQ1bJoiScMDWEUc2qXCYIDVng+K6f1
m45yP8yequzSQfXd0Qog363pbQIztDyw2Z368JnhooAZrjSw6Y+zdI5N7scyPVFv2YdwooeB4KCz
Gpb6JrsvVDKfDUb3pgZrfe0buxgx8LSIHf94CeqRB7+Xjo0+UgyVa5c0JGRsjpOgtP+3IYzlN2Yv
ojk4oFO2k98R36AAiUKVhhXWr0xIrttvq2K6d+T1JDDcBSvltExW1RlqSqA0eicM8EcDYXbuxcqm
+gXWxkqWdUtlWCiL8O335ijOpkPIqGch39e7QvEycFV4ywjsLqF0B9lRRsdrk//zr9kQHninhhex
Vfx9e/6D26Qlin81S3Jn+tRIwYwYIk7K8iUtGr56+OhncL1utIj3Id6YZpfjr43SthJhQUZpv7W0
NcLqQq7PISkA407J6xXzrSTwvv/50TDSVCuGDxocTMovUasvfSThpeo+viCLj/TyVIJ5BsRtF0Zz
VwnAPVCLa3OV3hSckJT5GgIvQWAf6U4DpyX6GHCKzJ/8UaHSOGt5xTUSNolihiqTq706Q2a/idUi
uWs/od2+oVaOp+enoG7oozACyYv+KkRrC1MiKQXiY/TG0VQodTOXAQgc2EBIq9gAjf0ie1dChIDI
FkJVzcqUeMHlEJd3kwR+Rhhsfuxm0jMDPlUKyROjh59g+aWOId11XBY5VT7FAzooNg7YXgZXp8vA
/Yw8XXYgsOLL4EBh2mjH2dVWk+EMErrpt0NPbCF+oJth7JBcmIHg9frQZgC2mpIiPGrXwW5lz3mf
BP2h6p/pHX4O1UAvXmPBZ1RTNuht4hGAQuQFFkBuboxLO+tsG7Vj8e29O8ccm0aLU0CSJV0l2ieQ
wi1z+WqMXjhTYNRLDTrkCjGVwU/2Y7GON97E8q3/w/jGGHzvrC9/z4Pe7EmLEf60TcBES1PR9tp4
keyenMqZFRLuBt4vjkNmKKS/nlG7S7YN6pqXOXlqPsbBS1T+/zC8TPzVAwTmPpIrLtfnv1gjpYe4
GRpyrszBsIuobpYIcBmAb7dQLk7gDJhqfANIGOiN0Bi/evMokLQgBAeXQvJBgj7ny9s4yMDvCdyf
u2SNBQaI3dNtg2m2hxhCYVVw43vYzHomuBeTNUwQoiIwuUVJyYTn3uGJE9JNB3EKvzl8oiKSmxG1
+pcEIGIznZAUQZuGoSHrXlFXoJLr8klcwJ/rvD1oQ6pjqqEmg4PFJzlmrF8TOW6asudBGKp4adyx
wW+TTELt1vsFYV4B0x6dlRNXCVQGnKE1N68Y4ZgvsCJeS1kvTdd27WxlrBgsCWG6XGCpKYT/kEfw
CVRTFCYrj4jeksoWMzGYNoLP/LBDKN7uPP93NAF4AwiUXrV5yICjXIkNwNJeKs+JOwRYeRoZjkgw
xIJRIymT5X06wCNnI6neyalGOIzTZbB7y+kaFfvmVJkAj1AZ9tKa4TJnXf3hOkJ0Dev9s3k7nSpL
jA76dAJcU3L56msKkBzL3rTo1HIogx8XQCbquWoFzUCtogPy83i22lh2Z1lQjt03z8nz9Gphej1P
Jrw0dDLMsW0GHS0Z8qp7tMY58PxXgcassUODTJkpm/mDsRcEawnInTKKsEcffJK7SWXRvyFXGILL
IPFz00l1Y07NYTpkFq040VbrGmW0pe0yzEp3JgDh83Kgo+QAzAKA565Ur2i/uLi4hLX7UM2ncALr
O5D98CArWyZkqQQ6eGOnNIgNFiBdBPlWssNbtfh+U9liFIyPY1VQ0PopU6Xoiw0qgZbCzkgcEMsB
3lo4z8IuEt3fi/EuTcTmx1c+9EymsWunzxqyTR+Kv6jUPVSVmq8sBqSxxZYALbqz3rbGZaY1RaFW
XJdnxDqtciVgwp64MmtBQ0DXSb4v49zytyNrmz6pqtB50W8UMwTfcvEVsqNjQGn7re5CiEIvysCm
rN4BtKIeHuB10U4nela5HNOQUtgMDPnzWCsOuyg5yhQGBSwGP0NZSg97jbs6sMVPZCm3PdKPwqo0
/lGl7UbyGyFEERKFNcN1XTonrbA5bb6nS8iYS3vp4RxEbsazE2IDT4HVmSTGDMbCTcwr8TVnVzmg
bvYJnoGjtoUkn6RRFvBcni9yui9ridm3zHcTd4KXPpst3HHnm8Yatt9CyVJK+NhguYnzDnZpPlkI
2WUCmuIoROvRVinw9r7LV3ywnQqG2iLLlDy9yaX5b5QiUosizfSVALaG/XrZwQX0BOFQKsEkrN0j
2iOTp88bWYfzvMlrIDBtJr2nk7LpmvKUFyZsi8pn423PvxAHdj9ybmo15WEWzMMrbbuQ3lG/oyv7
TQhRCznE736uo83YBn7wdnp/ejv/aVLUJOYNBH/zWGT5jwYH5dwdpfumrUpdR64zYTCcPnmk1c6I
nMepY7BQhJZneAve84oE7nXsDHg2/AUiXNXOJVUQEFOHXB1RjO9BH33tvacVI4+RKJ1jwNUfJYf5
W4w3v3jfrK8U1aauoyzI7O7a7xbm9Sv6Q9TlvKx1fjklNOzJpsObN7PjG7citw0N1D2oMOewd3Rh
6wJKMoArAGdrpg70P1R1+yJnjdpW+FxfN+b7bezQXXSY+HtbdtWB3VbPJSzehcISfUGwgTo8BGJ/
3eX5GXd4QUM8YYFn8MV+FQT7q5rvU8Cp6EhuNElJyJOHsZ6Q960cQIZeFzNS8F0LJAtBtp3yfOIQ
zsyyrMFXB4zLlc0Nppu8/8bgmTa8H5ejzxuTK/u6TICc7avgCpgiQ/e/Nmd9JQGeGPdwNSrv400Z
PuVGo0aiNlclzqDw7Rl4WFk+QuC/N+H3/v7rW4QBdpY2PlUY+rEw0JCCHHOt5/qgWgkZ3XESvUg4
K1NA6+4txghnM9u0MkcnC70+7lwCfAhb2zOKMYmd0wL6QaMcaLQ0KalTA92ELk6b7dHdaPTQJ+dk
H9Bagd6sRmTaICp0HcqfNFJmt77DrSCnubBkwAB0eAfYLSD6k+yDgEJjjb6QNYqVChrAI7A/Uybt
Sliijkb49UB10/Lc5vGvqjs71f2bu08p8s9exmhNMWrGwHXjDEsFuLCe85prATY2sQol4usa1GYY
Mowkd8C8pqtExopFKECk+abrOdFZwoZ0YUMMk2WPxJQS/DPfM2fqIH9gRKKRTymFAD3Xe9P2lJ15
FtcYLEWX+qCrTRM891oBUkbLg0o1CEyEwyVmjcftCcT1p/NF4sXKFJ8B67PwKE/DjkW14L/W5esy
BsPI5zz9cqL/mG82eSn//A6FgbP/WP8ds8MIptHmz5pFtS41UL5qfB0WxMXt+Mipd5lGmem4Ycy8
WgBez/MvB5UeOyPHQEgdtBJ4peetwEnRd78DUThZXHe6hQpMR0AtxTwVawT2RehpSeFUGRIG03tM
/1zr/PCWw2cyFB4rUW7iE97B617km8YXvjZB5IaKC68f10m/ybhxpnC+XlZzYTE/WOEuRM63omj2
jgtxnXRtebBakA/7k72Xu2tmC8J4emztOwFV++YI7zcb/v6K5vaEXK9QBE+qsGmnLbkXlgcA5I5W
zRNmMzFYoEf93JFst4eNPdAwLq/qvBEI1J4Pktvv8i5CLLuOZmUWnvvazo+GxsEprOawVqah+cni
xkHFKtjC2LxbYjM+eiT1AsiI5a53BJ0+mjO5lBZbbf57P8f8EGq9fgEkgz2bj5SM3uwE+4XfqVYA
hFYAD9Z1kV26tDpq2O/LY5LRIEd1rW9dLQPeduaK3BdUd3Dez3IwVRZzQUAB2H9hioLtZw97Zt4N
XKkMSrLRRi1pE3sloOJ02HfichuXIsAq4dHT+oT49pSeMfjwCKZjo87wmqh9f8N+xxajqYimLtPQ
3qltVBhN4MRzfAFOwc55bi2ZYG4Rozt7aJfY4AnH0LGBEd6j2gYzDrMiG2NxbdCpkoc9swIllkis
ObPxY+g4/+lWcNjfpvJEe6Sgyb4yEotr+A47mHpLo4J5N/msV9owUBEJUgc+dmB2Og6D6iLpL2FN
8ypkMiRZH/zeCiOIlAxFD7m2rM0LbpesgSQrEPkkp8cL5Gy+8ZmgSt1x6Yx0T/HSdgh8eUUb/Xbc
Accf7+3fl9gGH/XzZZuMTCuEkp5MYTRnRvd6RSDREUInmAhOXcH+No6Lbgm3gM4OyihU8yYDNKl3
35N8ozCe3PSHlvMVEMU5cm3RKeoBj9sHZ/i9/CIqoN1SW0Oo+6/FX7wEKcgZmn6zLeOJbZJWggS5
UDK4JE82B3zRYsuleDHEkVzNWVzLUxV/+VxQxVjMMRoZjb2zVLDl++DcqTIQ8szK8IN1OfNFwTeb
toZxRbUSkWC0Sy2eC5b8aaMug2ygDJAIQbxGcoRVdk/m1nZPPa6ztytQhQHWxvFrb2a8LulbtDXe
KX7hsJF2u8QvtfC15+0UdmL0zdf8+jzV7t8rFtKvqxoN8TNoSXoA7gkKvsauXmo1wwfERrefNRGf
VdJtLUfnqJet9MQ/a+obtVU567PJfFwMBgv/zAjwMt+NS7sGJey/NOihAdqvYM2BdQXOvDYgxnDZ
7ceMJ1u/7GITa4iSXMiQ52l0eg1PrY+58PBahpcvGaFNd/907dmT2eU7urB8kHihT/BaIhcm60DY
CCamV3Of24y7pQKhooLT3G0Ot5ze/AWG2kLvSnnW7nD+e5z370LAVyeidqenPQn8SkiH3hqpMI+m
hDSPSoy8i6Xvn1gct8hRrQn3omRn5riQy1BdR8acKureWfjqc+qGgQJF6iGuUpeurVT/dTjWq1jv
oQ6jxE2lQhIKBXorDFzP52fJ2m8lnDYGaZHWaP3y30GMo+GtlNqjgeMtig/udfQtUlKKi6rntbsA
Lv4Y3i/VPFG3DV6tac9U0Y2Hre5aqltpmDuNxI8WiWbJAmViHhrFvaUULU8w/vtqMwXjAdN4dsqt
bkmj4D0n/ASUoS+/peIA0G0MhFnuhohelhxO3EBjF30pJpEeKnVPahof1dJug41mB62GgfazZyMm
KDHm0wH55mHUNEbjp0KJyCJJpowPLRnY4ayy9L/ZmUISww5WtS0vs0jF0nOnhIUcZUFMyalk6sYp
pHu4NPzUvqdOzUcrs82p43iMfRmxZyew1AiAXu+nvtCJoqsOh8xLpi7GMwVMpYct3cOBaisWd0rG
UN3GveCXs5MvkrYDAHLAPqAyfJLDg2sFB/v1f6ld75/VM/RbdO5lPmOzQl1TotszwLky0gllakl0
dRRkp6/aoHGZMS548o8sxoE4TNvIdcq7x49EkNYODHty4f9wd4nrYzjFM02hW/KPEb1AcjJn+39s
BYmqsm/r/kGdzq6ktYYZFgkwFdP4AOdWOcKV2Jp2DAvAd86cbWB9dbDh3vjGF05x4Xo+Rf0Wm3vA
0ox1wRh4OIz0tCwc+EQ97D8FbIi05Yr+3SfIpXy8MK/iwAd6I8pT3+2OfVCctHC/Qg1DA8OFfoes
dYZoSHsfs7f0Vsoiw8NMxvDfug4bDAbjxxYPLuaHiZ6zYUrAJLvNYrqB6DfSy0BRD658j6FuLqio
hUFPneL/7GxgUSjor5Jgw7iTR+nRSdNwHStTc1G7ePw72AtlrpR5eUbg5tZCa/4433kYgx1wkxwV
luql5K5HSrzAtvQPrTLzbvhw4/BkP0z4VZooY4NvbWFc/77eDPuqx4lEoZOJKOlU4/4ONVUkPGqe
EUe5Ct0cR9QcaaKDaBra8r3cTu2o5kiaF5k+RlTsV+Wm9AmCvZbxUWcHy0gd2EJ1AN8bieRDDbiZ
HnBEA73DoQHH9TC3CKEBF9DzZpvVEibfVoPvAa+jNw83q1xirm32a0djJkC5mwSKZ9q68AnB5cPk
IfsJJTlQIH7S2hdY9JdAidfEIi8rOsZr2s5FRzf1LyYbm0d00AS2oqWgnFnBeXmpN7IbQuaco0bi
1pG2snnWNSLr+W9HAl6yJu/zMmcHI9vBPk6lvjnOra2U/3Mw6Wvv8jtyAjv1CjtEpkTc/W6i4ruk
chnI6vRkQCql2RecIEsLwrP1SOFN8fFQI9+66cQCP3x0ftPDaHJsJSBsIfunxDjWB21V1VH52haO
bYwITxxWUPo0+a5OJgFm4QsOOAlMWsndSTDlEZyCuCNg2OiaG3MzZgSVkaMxs4lQQkSZlm3fu+6y
quidEK7KhaEqb66e1PCflIuQ6WerdkbiU3y+E3XOp06m5Ls5ONtZq7oGCiK1hBGbOQ2rC0/YfIi4
pgrlFl6bnH36h7nIQpaCG+I12X1lyTLB3nrEbgazIPlug9uV//dV0nvK9zbBmO5+RE+nqTDCpFPt
RIZ5KwFG8aSs3/KmnwgsGFSnv0NNWis+96nu7O0o4SJ3V/bWXxBbZqNMsNgRmBNUuS6PvTVkLbWP
oIPc4UpzHqp84GTgZ8ccgARMUrn8UXZ/iluCBzDdQ1FWOvdZq7S3sXuy9u982NXH411zcJrtsUSW
aE+woylzwbQ+BDxg7hE0Oy05L0xaVJO6z7iblH3J/VI3ckfOb7n4jqfbLUfAONXiAYY5Q0slV8gp
svlXGZBMuzZWjNujIcrziC1e2GOiTNGJyQPdwOuU4JtA4oNHgQi3ur+e4d9Oc9jQv08zW3EBx4ip
D0IYXLZ7To7nGn+6/7mL300g1XK1wnWgV5WPIMOl1EujET6UIUH+gCNgDQVTBDlITbzicCxiKKg1
VADDQGSef0LOe3dErPwhLbZbUDzKKdcrMx04+QKJYKETmUh8VY5zyJzCYMum/S/4b6jud/h/k79r
lc5qHzhl0rpLcwQrf/euR+d7YaJdouzPhcrm7t+Ye4KOax2RGLBbn1JYdvJMWVMQ3cFdJMyXmu61
zfAfzNILlocrM3PO+LjMThHkpV61qQ/xSSHd5hjIWjYubQTsL0h0ccj7p02NKk040LKKgBX005Bp
nD3JPNY7MF2d/qCoK2py5Adv+sqoNSvREo8e8L6/BpjFXUcG1HZlOSCWVS9nZH5vXZm8atv9T27/
vA4kCkGrnX08NE2k90ki7COUk1RyMPzeZFX+K9XkHgTd25sEJ7rlN0duBg9x89S3Tbtylf8X4cbW
c47MZW8RcQwj6PeXHk1yAkkmOzWgUxKWO5tfengvlDperWU5zwUiNQn5MhGxKX36VKbEvWVyaF08
PRNHzjt5wjOxDIxyiH+ETox6czAbdFT/3LnYHrPvm7QcNXywAqn6hu50zCa/6HITKpwC1WWvxrkO
rcb3OBoH2l0bIrvE3SsSR5l5HFGJ7vFlsXy8SptP1+lUHAoOKRq20wavE95BHKFrwt3YFsMx6IcC
fwyDTlL+5GQh1VQ7Q0qi+VOctGxGx9S2+/7vSocULeCO27wtPEpkmZqMktwpT8flnj/1E4puxNOT
qEzshwhZBVIZvaUosR20HeHPiH0/fZlpdE35PQuWVF23NAME49UBlzXAjjtupqf58wmm8AcRaJf5
CUBLXrLT6b45/5xeYbzD/BJctgzcvvReAZM7xJVS8JYfokQ69UcVBpuRr+1psCUil62LWhaFGev7
z8xJWL8eK+e5gpT3hPoFIpleC/DLJcrCOkHHs7UrJRiWd+/aDphWvJKDunj3f9gwADdyOUr6jfhU
vWbDkKajWQ19Nakjf8tCxbYnMPHFnD22eycypQXIjqIZtb6OGPkJhtq/lme9DUZGD71KdHGJc5wZ
d1Fb0PyE7AnxrkX5GE1AeijlJlC6gk2519eipmctvMXUvBOJ0WchylReeEuH7y5dTYl1dI/VJQq0
3ApDHorzLMD/rBtXQjdum+FUbGrmPIRQ65raWZIEyfoCxLI07wkLR4maVVeNSYfuQRjIfnst+v6d
Qa7cqEWN2gFdvrbs6NlPAoLBb6sm60er56ggDRFatghQfVwOXb5Px5JPId6G4agnEdoynDMbOXa9
fCB0v41MrVy9urLO4q/JKdlWysHIWyTk+WCtLj7RWyzyRG5vZdRbPAvvyezyJMdz2pEcfsVCqmcS
1/BSIg71Q+98SB0BvbceGcOpL8NvtX5oMb/I8Jm08LCtcVVGDHfzGwoerrjV1+ltBWDW+GBnyqmO
p3GleUFmq7uwPzMYwCn5J/ogQfsuM9I6Xw9GtSJAi+4HHg5IsXpAIvhbJPv3D9m0zJNQgfMwFAWQ
IIKEV0Kou/Hklh/s1n2bWdln213wtoTULY7zo9cnccfrfBgHC3rI9VGWi8Al+0xS0yWV2+iogCQ2
ZUrKTpLwSIhDFQJdCD4VlTRShW5/LP+Iej9NtxUsLX6zagapyl66S3TlaKcWa1TphoI5z62Ficbo
8YXkPhREDPx3a/B7fHmhcMc0KBAmd2HK6pE3msIOs+X0D1exezysbnlwDOx6m7RnxPYu1+taT2rJ
FUfyAtUh3LtObul8iEQPbvPvfFJNCkA9974/MUM85RYhkAegOM72p27dTv2B0ktxlqGjSDLoTZUN
neFGAzv1PHbmBB7Ey+NS/S3uJQpoxHM/fkFp1M4F4d3F3hYyYCciQ8cMCQ30GDVd+Wtw15WK8R3I
KsOajyULqw+XYSD/VEUsMyzTrdEbngBHYoNeG3fzb757aqHhAl6rGaDDqn0oVKjkStq32HOIHcH8
0Qrg/E1EteJiGt6oiTrBAff7h5qh6Jy9oN0LlHWQpuNYXf2zqIzszRu1/sQzxczqcC9rqkGyZL0m
dk6h/2yIg+2qZicG6GmfbR4eSSG8R/h/z988xohJlFQS6g+uVJSumj8BaTmSMVpqFyADPvo5k9b5
Mx6QPsQxYl3yTaMb5wkfL+ou2AWxl/OXrqvLAw/uEpE04ex1u7VBoeW2PcZBRaEpUre9eVApUK/c
ZNBg1SRlPSUfyg6DS4OL/cetNgzrgw2H928pavo8nXstSPexGnMYlDK7d7JcCTC3JnbeeTxuiaxC
2J90kQSQgN75g9awQbU4GHFrRoArMv8OTExP6jHKnFsvlQ7LOTrJDZqIeE4KR8+CGPfeczMw1laI
gIadyj55QqE/bV4PYUd6BkZzwrDsud/bK9rIE0FhJPgqlhLkp7iC2uTfE3ULYLVSBYcqKJ2RJ4i1
JDWmBI3rhNOBpSRQsSCeuFIfbWWALlSLrC9rsIAgvu3KMBP9OQnmu86nBIhBkHtEAlKoZk5EKFqk
jR2rtoPJb+ZqLLhn1FgwVkjuHm6voxGySvbVzVpkxLEj7MofozDV+LeuVebOFSL+8jS30MCeMIPk
ZE4mZ5tyxNIvjykJaw7MNZRPiO+RDYsE7m+dqZFguAmkxTxHR98mdjurTKno3EAZsoyv+vidLVMI
GP3V1zWbI2424ob59MnMc7Ie/hTzu1xOMO41/dhKMruKQbrGN26PufOxnFgEtKIWIwuyxSs024gf
T1GKziQS3AACR3+cHe30u8QmVKF3aOgeeFGxD0vGhqtiDAsTP+WGWLzPwxnzWKFr8ci8X4qFKYr/
kesZhgtBDhLx6g7jG6ISWfkYrpvgVUyOPJiIBp9jzr0s4dctLWouBJBwdNobk4+eejb4kLxc210w
M1sMzFUqLrNd40hboMoJEWO0mnxQy+Bh55ZFkLQ3m7G2cxVoetwzqB+t22r2S9+sdlsWIwGR2Cgx
PtYHjmDjLx0plDXhgzXLe1yo7drwHkdIJ+YpfeE3ybOwt6p/kRFocW/s+zfZuZz467IwSJ4798qp
gP9pFBFco4mLXWcfuijZ6c84xgLX89MzUq0CE/hwMJGyDfKyqM00S6BOGkCPVZrzLhksBnLtUAPu
DSGzocpMGcHvXTG1rHRTMkrQIAnZJxvA4zJjOWxStPsGOqpG1Rf3VQa7SB2hCnxkJD9OTn/a6N5S
RjPW8hv2JHkROy43COxm3X153+D5FDCcxlwBvDap4DrcZGMaeBnMtJbzBET2RBlOUdDcscpFc3WA
7TbvvUsW4E7HdLwMpI3Xs8RodVH974XCRYGKbFE77oh4afOO1GWSauZIhR3NDP+hb9l9s0xjACMY
6ATCzxzoh5COcOypRSmEpnnwI2fhDFO8Gy9K4ygmIfh7B7ykb8hqIsiGrjPUWiLD9pgfTulM35QJ
QVe9wi5p+5kh8A4Xqxdn4wSlhHVHUeFZzsuzebsyTSLmY2FGu7Kg6QoaxL0ymMdQuF/lTxhqx4EM
19Cu+SPM3sZsDc/fzg9MjXba6R0jnM4m7NVtFKVlOLwoUm2fr2Abe75UVOvG/kXrlfUUIRAj1ssm
uBgDgjdWBYwX+LbFgNesJt2tc+6fEW5u0WYT9glWcNY1wpfMhQELVeJ3AVRclPDgZdEAJ9ejEHc/
hQh2WG0tEokNQJaw9jKswVX14B+qttLnNbNFCDLZJNoW9HfFTEB7J47CLFzrW6gfX8inPrES9ufj
nqD9+oCtCeasbqiTkFWMrg4ZScJdLV8fVl+O1mDorbpO3Z1nziyVvl5H4xBknGLo84pvYbOHW/hO
K3mhHFvF04GiAwpctRGDOU/fIlTNcxsLTErXYCC40hmOe2jJChcrZXUapeupu5PZbgrVpgdXNcG6
1v/fRZQycoPt2llTzWUSXfAKhzsqlM2zgyi1oSU/Ubsygl7mp4wG4SyuVy/wOCI1b9xn6D+Wwa1+
QV8GIiRM49t5LI43W9rXLfqz3zTpm5AVzBar7Shb4F/k4JBhqRBKqe8PTHhToyC42SQvMtI+SChj
77wu/2ZRkDkS3HR8WLFxKiodVclCAN6cWNQffq7zEzIxfndDh5WJ9Uv0iqp5lEZMJap82Hmz3UDD
ScxB+0nCWLaEtkVtkT87owI6NfYWS1HF7UsCcG3hvQ5YCnegchUXNWFXsm+anVp0rr4m+uycmt2i
RIsU8sqUA4+TXRg4oKH0yqRO3/mKTNdcC1SjhMBmFleJkA7OaYiRVuc6LQqqluJoTGaKxS9AA9JX
UfFf2r+AiDxwto325mfc44ErVNcqkOfyA9xFNL106MKJ9jpb3Y+18DhqUjXE5TKw8Ib2LiX6OO8f
1pFUITXB1PIEENtr+X8pJDr87CPqSoVd6QXFNpcca0/9zDLQNPwkCAaPBFAO7tcnrfK+QN6I+Kng
zX+GTO1Wz18eqx14Ug8PWDufCbw9daMEp2gr9KWG/+BhfcQ2E24o40JtFITCHlhKjmEOUHsCQ2qU
GLONGqkpQszGKJaiKHgPv6rBltt5/qE8C4l0UqSjXg4lcgQQeLtZL/kMcLG4sF427VWdQyma0xJd
R1PIDjoG+osTWLvZRmCh/XWt8j8D87kNng1MBJn2YSq/HrrNYyc7pZGn8zaAUX0eFwaw3BsIXxdB
6UA3qO8nc6y6ezBLIX465+T8FYWcmgE9U3P64LEF5NG0+rrwja5N7RI3T0bu3vEaJcaYxqMJTUFv
aui69qSISz1n8CrMruWANbimgjox8xFEmYhkEiT6OQwcyCVPV8Cfq++1s2h8R6z2qLh8KzIOtel+
j3MqQKTL0LpCNEdWtePBZxZ8ZnVGhaR+3mGhYJN3q/V/GP9obezZBG3DwbAcjU2CaS6TwYn4qTi6
VFDzhnzhrH2AHQHtXPDNX/Jy+6aSurYx53BlzwPysonmPxtCEg4phEr0kt72Ut3aOhfWAaSUK8po
TckXA+y4hj8dD6nYnXoz/8L14p3rrULYWQmtfJPsmIsn/Pp2Q4S1uuxyeJRNzdakyLJ0A+MyV5Z7
PSuNm2TUda4mNCAtP3F0X2eDrl8+8PK/UxPzw+30UEeJ3GWTGJEqIZhlZQU4Bdcb6473b1StrcmX
1AcM3ZxZnKHp9/7hlVYUZqrSuEp+3vEIuHiw/iS7zqOThZ+BgUAyehmLU7SEHBE0eP0vt30wx8af
2zPR2+GnXonVwgrZHtG0pewPeC8ex4A6WSF7E4LpqomhhVTu9+O2Iwm9rKKzB/zl9D074+c6uYY3
qw5MvSCjqlTwvoJYjh35iSueKJtf15qnkr0dSu34IER59KsGmjHtmG+QIIuSGQx5jWaZQQJ2vcVi
/fpyKPNx5GjvujU5iWx/8vxRWhyqOjE867vXRycNydO1/GfXPMdo++iXpROIAS0D0Yspfp/5Vt8V
PZYpWHK7BmRtOlhsFsMAvhDi4sEHbHT+5DUq01IrztbmamRsLVxH4R7X/VCtMT5/9EQr4ScR0Zrs
xE+dyKLh5LixwhkB1B7WoKwenGBwFJ05EkHEA+hPsMsKttb1I6HIXp2fKGtq0MrytST7Vlm1/t3W
YQ5LboKjs7PQkKuN/X8ZcmX/d4CJQmE6M/fvTT6D0U8eyaaFEIpwb+q2CRXfdgNvlDZ914gwDQk/
fG8tRSMfvd1lD2k0spRzKw8xEcjzUnF08Ah6ujRrJ+fYrdlcETSZCaEqD5QITxOZrV0fNTqM/qqN
/faTnv/OYz/V+hwKxjXZKDnR38tgVKa/GDrACt2hib4FW++FlilILDafj6/s54B/eWtHeRBIvzmx
A8tYUj8/knRC5O6LGO0tYMi9qqgzZMspCMfkRc2R/+hCssujC4GN7KVWGSxA+O+oYQjg5mMp8kmu
FJH7DTKwS+iKBKOZGV62hCBzdWk8rGXPsMv7GySUaN/dQEm8aZ1JygeHR0tUvZ0uTJSZoM2TqYgM
k5Gze927nlrrQUBORdh1zl6GD3yzeSyIhICJp2YXCyDO9VoA/My/0VPkRVBjMnDX1kX+wNrhxK6c
r/vv3u++JQSLDcYRtDApHJzGRdXBCLtBcHW5SSl9j7CgCbA4mycX7s6xlk3Ms9XfVZjjQu2opbHc
3wbwYwa1ECI2Xfwi6YWfGYKWvIqOfkI79D55HIP47/habjxrj7HvMFWfAZM3HDWvbUuIl9Z9wlX3
r1SRD4cJnDWjNXUhSE0wcrEdMlczRH/Hq+fqJjqoOeRh0+IWQjvUa2oSj5GpdMbqXb4M7CeRrm8W
FrpUsfzbgawpNgGu+dfP70YnHOWJXz2vaye2/8vImNNV/E2doUvW5eU0eW99QXE0TKBDz10UoV1j
Q54G6XnTLPlTENQi2R7zbDQyz9UwTr9dOgMu/bIR/m18T+U0P5PHx7QiUMlzy2O2J0OvsFM5q8DF
PuVGucokihZjWfzMDViY+DAyeLITXzGsl0JHeFaAXWuHjFpt3b5On90VRYegyjjhj5MkOX1JwK+v
2/esrhhBk5Ajge7QyVf5N81dLIs6saP6Wogpg76zatWI413bmmhZqtJsuM12/VHgO0qG10rTQYeE
v2Blv4KQ8qUP+8ulOcatBKXxJFwaZadBhjYfNK8xY25JmZI4ycqc2SsdPQe6WqFfvD8eS5bdBd4p
x6+Ms4X82g5fIJIt8xayLTi1KPEwCrdUQ3ZNRBoQkDcHhhTgkqgljzMuffeKQY9PjQ61rDKu4tiZ
d6I4Q83b6DSZOkAuNgILMPm/dFjJ3OVbO2yxEzlW5D09N1+FXFnrrSIiiKPox1DVGxsnQXECjjNI
yrzGtMOxmvuEp3JPtRyk22vPCPDeK0Q+WaY9kJN6S8gXhzRd61tbGGVIBZx2f6lsevF834uVPkTR
pMhhbXt9A4ObNNsH80w+DtC/OIAj11Q/1rn04ddZcu6b7X5qPwG5/RB7K72syRP4aCj8uylbjtzu
TxALIRtIQGVc4bLnqwAHmtBwzHGRljZ+Yf/gO5TWjSqFdIFyg3p0YS34LDw5Q61A1y6MJzPAOzVo
IF5xD+SaRGiutuVaa5kBZToG0LSTcUC8agUV7oWGSuWl8oSqM6mSgOR0JwTEkQrtYxnx7rDEQqvm
6gb3DWQ9jy1DhF5l9LWZBqtNgB21YFWd6TL2toCDjkjLz0i2sY1u/PegSemVKLqyWbQM0U7W+Vp3
c7w/8UkdTcXa29qAPiuUtQg2XrgiHfVrDdtDZlXvZyZMR//2P89giOaxJR44UQIjbkhgEWGpTN+F
SAkVxCIsoLLLEw29tOR+NgW6A2OMnEqexZtYkCKQ8iE3PJmD09ijd/7oJE9+AhPNQoRSfX0V0MhJ
3ioRbGVGDEbmHgB1UEVeq91mN6kCKX650mWN7VZkJxftzakNxBT+IeVd36//llLggqiH3IuiWOb0
KCBC/wOL09XoPv/HEIAUIg+FDju5AzaMQ0GXhJJ86zp4Wgh0FbTgcEU7p7gro3//KGpnMAFATJ8r
zNgQ+F+7TIh4PN5+bVTCJ13xvD8Mx1RHu0I2R0nb2KxApdPo6XOpiYIyWANiNVryV5Qo/n8lYX10
0bE5LZSACxV4EOQGv5RLF6HwDfn7/5i1zKihKfeVqx/qr5fYUQjj8X4DZfEr591J1YynooTojlDn
uOXYAWqgDp8tWW3DQ87vlleCYwimx140XhdEgCT6tlihxJ4SU9ki3ATOUWtejmiE3FufMBASLPe6
ZUSpm4NXxO1dupnRs4Z/B/YnAGwe+x4GCDWzCIAo8dp48sF3RY2SjspNzI/IxEBXh/ylUOEjHO8q
Vokh9w3MlxCjR+TwAhm1pkYn+baLrgU1K+bTsracbLiF23TQncOgxDJOFvIbGt9V4OY24NpVl8x3
g2Vd4A9jGBOts/Q4WHsz+fyO48nqxJMtc11FYww81l1evxQ4zMmtGQpYIAb9HHLgWChB/NgD3OUE
uIcDgoIacFHC3k7Bx94qUjQpKVT/8wyd7uxB1nc7xAeFM9wEq9sZkzZba8BTpIcrzOq7YaTJEc4k
a4lGO+ZzZgX0Pl78JxnNnUIHvpZnmjavOnkBESzil/rc9gjTiQ62PRwTvlzrFB49Uf+4KFByZnrF
TUfCGMN6C+c1aMM6D3p2t+LZ57ilic7MJt+0Y9RbU4dixZ7Cd4YgASgq3Sg51wbfhSTmcvS3Oajh
Le1Tcj5ohIqvteUf7d9n49pSNOvt6IvZBipVugxiYTEJUOhI6XH2Vxdx201pwn2rGxe3uMAp/y66
lLBrTx9lZ63Qc04diPwwuMM/wcN18Lc131wgundclrQ3n8CUOE7mP7O2umKPp72jH0PaDnork4+N
OvTvspaK2mWVOQm6uWwNorfJbkCL7AIcRGmWFPi1tKxN2f9EBMUdKmrp8piMhlNQO4OMUoFciFGi
PzOuzPIyCho5qOtkCJk0bSIy2dTgvJHsIfuofnDDw0XBNcKuqmHtxxXBSKuh4hijiwzjBCY8evrZ
ICtoy80B1+UpYLp9YsqHqelF+In5QW0UdZq0QwF7ShjorSKYC5LSamau+D2fkdXifduWJvbdJsIu
7zpM8A5HfvgH3Deg8zTTbTSgZZnTAa+scKA6IUKAjUN4BOdXQPEmu/3r58bxfscuq0c8DHXniBDn
eV0izGtBoHsICVOZhRcL6yLXChT9yVh3P8F+JRTyXb5q+I8N72rmEhZgWKWrwkdJUsrRzV27uXNF
JphPCtBk3IgEfmO3uWccSzqmu3zOx3CaZrwCgmD2qE9vTCt4plyFkC13knYAtH59lr7V34ytEurw
mJXwhf7ook5IFSSsr3JWS8NKx73qd6F/wIdYQYNsaqIpQegS8FM6Y9pUNO4J4d0586VZirZSRGuF
dYSe0e2byFDDcBO6ZmRz1R8Pe1Dy80sWXI8uhVBJO7AcLQ32ZX2p/Uyf/5K+1YvfGQbcEawxIHrw
MAdvjb9pOYSDTeCYlFUjS/bSf/tI+9w7zS8i4VLPZpHywwt77PCulHsRYPU8YwR19yiu8JJp+un5
+iF/IV5R41vHK+n3QE70T4owhNGqE0QHzvFtQD6bO+nEiLkS3/3+lQTeBxyKHC+/JYvaDs7UyjZX
vFO9l6++XdD70X9lHdHu9wRt1o2lrRzpyGqc5wRDmmVOMrXGS2sJV/bxf77fnN0WbtuoP1YyMSwl
9wX+ijPop5VtZGjBjonPZTVXCwMpg8Wv3ncnRbu4SdKlbqSGgy6y4pWbT59pDk1MqsMAGA7i9Wpc
xykInp2LSH3V/Cz9MIuvMuMq8q1spbZ46JWuTddZdsD0l7i3l2w4rFwBPXbGs0ctuIzS0e7EtoLT
NfVMPvFJ07txVz11BQ3gAnx6F8lxUqmoEQcfQblAk7HFoVfAkf4Ux1zUw+dJMgHbhK0Ns00+Gu0c
A/tGMKAqHbj9VWA5vYw1hjQ/9ox1mavG6V11G68wSUq0jsiT8416lYON6M83SR2yqbxdhu6mSrs+
hQkEnvLuRgY/PhC2imK7cmrY82CVzZrJZuisO70laNn4aA7XO/OHRv4AazSeH2f1LLHDMhiTJ/6q
+bw8ZEzckInjnmpDc4DGwZmTeG7XLXYnmcuCVJvRHSmvGK0uBYrubIKsMZvTIeFJpdvC0V42xqBk
QstYWl4xBJNEriNjPbXv9oJLqr6HLR4cFPMqawzhRTwQnftrFYS0nNdFriCY4Hl5jIjogRHCTgtj
AtW7PQRIk+ogBNuMf29xaUTflDvDgj6Lt19dV9fTS8NyLhuiuXkvf3MR/Uy7hhFyuAnPmEzO+wGp
4ie2jIX0P7fttxhZPewx+VQlKJrnwb/w7JR1hpn+IWryF5OAVUZqYBK7qY2MZfW5TkHxCG+DH1cC
NtCaAWLhvgVPDsUpxjP/tasINSRm/GR3y1BXgwvZNLmt6O38hyVR2QYlvnqTpgKUB6WB2mNPZPWl
5pVIqlAxBOxqrl7p2JyH/f51ekAyeoBrKaQik6nLPJgu6GjIfbVt+9q7aMgKwjIDDUsFVn4ABSdu
rVRpgx0Oq8v3awTSwKKZVVdvQUsQzTuphcxadh+uZ88gH/MqYrphbfnutUWtD/QbW6ziBUvkGeMo
J3Xqu3FaWsYV6HzfCuBrNP4toMTQTO2qQk8dUa0iXUOCUcIBcQz4W4kkQeM9ojdEPoY6NUoGUAMm
mul9LmvgYBUzsteS7aEUgPrW3uHJ2qwQe9EdiukHiJB/V1sQHo8woZ49N6ThycbLwo/7fursOuAv
bTmzkAJRgO7CBxq9MtJiqN6ElQQtdV5qYUC0BTNj8Hmk8C+aSERz23iJCIPzHpt2i5fm7Ryu+uSG
WvbB/94uInB4iIsyHMnNS+3f0tEoAzCRPM+2FQmI0dVirvXC9kcSFCs2TFHz8FsLdIVtFcL2n9Mn
3eQeVuNKjyoZBu0kwm0UIMDUr6vf3XBCY7RsG1hU1jZkn8kYAVtLhpKRJEsXa0H/i/+DBx5rv69m
rGRCyM3xIS0kct9czc+wsLJ8EG9AjdnRoBnbyR/KBIo9EyYBUpBIhf5wraff8Q6nZ1AKg1UfgV7E
eZrLwRjRo8sZQs30zDFe1XEZ2shGTnJ8KxU0mWEPLS+FaUKkRAcxWx4NItPVIcouiOAE8dlGwTAr
gGUrvQLkXuuOjpQ4VfNdCeCHa2EZVEN31URXoyCdEkVQQwlQBenzDe4wrk/g+5eqiMeQeFd0/xz7
lOdgfd8o0cidP5sA7R7SbjDlSv4CKxE7SGvPREJbqF7yv0L/K9fkz3+rcip100yolz+6Gbv52jlM
IiMv1DKKVVImP63GzOVhg9JPOIstUAsH/KtolTFbbHLEcoASEO26PyQJaXSTTzzr4HysqBd14TZA
aftpgI+0nbus50OZREXoMRDZmBRXZ4y7ESpzeMW2gL79c7rDobrQo1liqTwQI5KlwAE59mhxKkgO
+s9V8oDL46CdoSGxikoOARKrFslKwyVnJsznePrDqmMI3N2QQrInSH96Vpx6HK1s2HbfnIdIT/Uy
mfYifAZecpBtkxfJpZwuxcprBVI8ctvQev95kNJEHdyhyGJy6jzI2/I6VpvF4rRPtlTc/RC9NNNH
/eox8aD4B2SfHQmaCYghpZLbYtVqVYVg3p37WFqx4FPLEh2DkiizBZ1RQo6i2c/RJdTOl2tn2GFa
VP+eQOlIGju0mywAPqPagr19yusTh/RP+TJ5UvzHMhavZthQnX4vWwXy996PsEUbiSmVc5t0BgEt
Q96RrcSuUlwvlzmJ1Mj1Rfmv+fzHr3uZOP8I1ntobrAL4vvRJoDCE0+Zl82X09GmeGlqGNuzwpN0
giS8G0KeTfc1PtmosXlgtJ2YFRgH6fkziMgC6eROfD/IAfVB7hhhX7fn5tKPOIflx0yJKB39wSrA
qrqVH5IEWLJ6BoObIwqZdG4kBSKazr4oU7xH0NrZeA+Jdy3NQJsZT3wTtvgEbtgxBetNVfHa7e0t
WBW2ezjcdeU0WrTu1d+yZnPhm9IO+aVrQGHzhYJqMcK5btCOm5yGc+PMklLOEMW+gPYFLDHAMzhL
mDmctFOqPpXDRd9DWqw3TA03RZJsPH8UvnGfREB68QwHFejXixL+8cPowdlS27R0jyQFGtGnHT+Z
HMPhrRcc47FdtNW2vRBfaIfisGHdebld4+IBaRAStcdxL1L5/CRHb5P1AWk5eTs1xvbDnOKrv9r4
fbZFadSzFqGRaPmxaRB2OgJhxEEfJzOXG1Eg2XQCd3BjKY5hzEEte0Qkjrdz1j+/1OFpVoJeWXTM
QCdoNQH77Ymqlp5STTutHfH4FpXYh6t2BD4auRvBkXPlj7KNIxZi/QLyBeXIOMJ4EAR66q1dnExV
ucRx4IVerlcZfrk/ClbhrtX9BFpbD3RkZbqtQ2GuIusJWa5BODrR/3UC3xm16UTBLIJ7KfYEVArR
M687shlmRGnG5Dn12073Zc36eMx3Be5+w/Row+A35qu+rRxp0tPGNhoQQc9cm1q1G4N2HX6qD4Rw
LpdXbRnX4HnFQuVxDoi6m8A/MRe+AI5za4p+Z9mZBkOOTdJ97Hl3lRhCV7tF+t5jZM0YWPl67ncG
yi2DoeRJIvb8FzzZ9dgbxTO2IggrgHlBIwXEcmEHcNZfErDW48Iz08GgN7nPKPb/9TnQqRiuy7ss
yZ22CHjugwgUH+A3LNQyYf2VBPpTgIG0j6oi8veY8WcTTolm3/UYGPthS1cQrWi/hbD+9Tn5Uq3H
wdGceqW3hJyB62eBKzB+K5abZiuiQOq+kMt6sWhGDeqUG/R1zzguudc8w7TOCpssME2Q2VcnhDCX
e1hEcvVXwmjp2ssVW/lGCCXEb0cTxxvFyvdJZiU1sQoKVCi0NsHpvAbOn551UsN6IDwwXXoswu6s
AoPz5bUkgKNT9wjlz6vhZ/8lJx90fbnnr4EITK4KknH0raPfjiQTxDW2Eh65NVz6yI9iy+KyFtGA
RMjduO7WhZjrJsiKSDyinTsgMFoB4h5A8NMZ2SUE6gUZCOL1T7JQo5MkG1LaHxbApXF8RIv+fXY8
eev9kpZbaMCkN4urKhoJJv+OZIITiVbGaRGpA/cotS+rkPeMs4S+P5dQoMM2NnTn8ymlfHCfNhgQ
az02Tztv0qOx0LzzyVNsIvVO+42izZ+S+2uCz8hpgt+m5hPdjuiIuVio4JO6w1KlfqoZQpG0zlxi
QcCiF5q2loFRfnMn0RLcMBykM9F0KhrpB1Jitv92Eop4WgBfBA/7bA9E9+aGyJ1tdRdl3NzKjLlv
GlPEjjjCnv6Xi84wsQmD/n+RQiJEyhwsNPhXFRIPHbH6GUBOrXoPQgMBJsEzlL1HIPpHquYM9CD9
wSADlmVRb/omq9zzhNDIkGOTY3d90vEehb7N9t7dT2uCroCzL8V5VUtT6laIEgAoTMyaM4KaHIYq
IsICiM4NrKykDvfTSOjEHJrZ/QBBy6vS2n8sx9+rc1k/5CrTnZarpl4ukxKg2pjCbX16VpnRdypk
JfBFEC4GRwY1VRMM0gmguvDZ46baLjL1VwIDQx4ElYgS77X+sQnt5h4OjGge9eGM1F4NuknAvyL1
pvGfhvlCe02VQ+8I4UAUQRfZ8wexw25XtZo66B0bBP8UArfMvYuzvh0OsvVZpNp0nr8+PDrNm1Cu
Eyf0ZoJEYgLQIzYpRtH1NYByLxrq7Pq151EM6gZhveKYLx7YuicnHrBQZPSXp2BuPBjnknyoxzVX
y9cKaeKz5V7SGVV2B/AQptR3HrQzMCFLPZXuBYLkPePMhavW7gD260tXMycFKVdGS3ocQ46qP8Op
vL+V4nsDmpj3ujXM4QVEikr8fyTLlp2zcSCDy6FI2m+phwThYDBiGmviOH0HYYXtFv4VRHJbO0kx
SoOx+O0rLTMvoQYinaoFXfrMXAsmMoYCi/D0fX0yYbgWXd5JaH+m9UJTbcuTkku3aYRo4TIO4IFL
7kfIosIiBzQf0Hxf2lmsKec1Ak9VXz0rOMT+4PN1biX8eJ7ddjO1gR9c5kTzcJcmJQ7KhSMxGreL
8EbGUWLviQV6b/AusmjpmJd+qlkC6C6FXnRUYGm9E42ypFqwkJE03ZWSRyN75DCch8r9K2CKlvkV
plwkwFwPXa/gxxr33ME+Su9jdsCRYJzCfIUxTECRMegTq1XUVu5Qz8Ol774GlpnQPceGEJ8slnwS
UHlIY2Oxvu+Uo5GpKVnAvf4cjsmSX7iMe2SHBbUFtZLuTgvVhN57GjfJP9AMxH0QdiQkgk8Ir1L0
uoZxXWrSzZeNQiCjfNz6vxoC+TT4itPgKlIGVLZBzUY6gsmt7pZirWA5nBOPMUyb9ZlVgcJXXGIm
BWTPDvE8oiOCZdP9eOqqFxPRdPP07LJUe7n7UG5KS1yG318oJsLEeD0hPo9MZh6dGSV32gPuQm/E
vqVpyqZIOXWwoNUMA/hoaD68mDpCcQ483kNGZu1oYnl+EpHxMgB16lRljEsG2WjVeyZs7nT9s6jM
BH5nLG3a8X2A3ojKjQ8RJqwvOGUQlqgiz4oFm3rBus0JCVu98O2ZzxaiK3MF+ZVZNGPsZ5Ha2HZF
EwptaeAOmKb9Y6XymygzPnOBIa0hrK1CtZaScjzvxfz0wR3PshiQZYKA/Ot8/ys+LQIsHFGUzwN2
h7qx+C1yNVgl49Nk7CREogriu12xX6DclkfJ8wt89HW7sI5TfGMYJk36G5xPS3w1Cy3EVaV5EZdC
wBNALDwCm0jPm9u29pE6RFk2v7RKdEubedozTIWeq24lrbGhgWKRe71scNJW6A9qUlonoXtykNa2
pNrYAzUZXGK2fv9NhVxe5VaJA4soL9awEm8Uin8gBfrRvQYFX0nyBrONKSmAT8739SOzyhw8RHHb
1gCPYd6d/8fetliU5CDb4UqDkIVqOD9xyGevbeEp+4ZK+IG7qMeDf1yKLrhOO8OX7h/L5941vB2h
qKaYSYWsxptc9Kok0UlBBwyO8Jtbv/P38UPy/uOxEROx6fcs0EL3enMp3vlwyrkvnsvdSijEZbsA
sP0rJ2rXdMadxNb0JHKkIVmMjXgFtGmT5KZXVOADwMoRAI2HtCldguFmn+kY/MtIC+MUAopJQ+wr
CEv20kpElGqKNDUR/xYNBAiVvJaNBs3DJn56yAniki24ot5hXMpXAiN/AK9eTIeeBd8Rm57QH1Gt
HrGIN9J9fpUFClo1ujjQnwPFLqShg2r0PY49FsRLIIq4MxOdsqwItX5MFx8j6x6oQZUIQokqzDHr
obqzPXm1woBklUALfZRMlHQE/Jg/vrFgWSmJM0Mxiv7gjHKI6Qr43iCd6+CIZvlEHGMY2jBbP+YU
NjUfCxvMfJoNHcM5wq1lvQ1sMWkQRsrxTNeggHyDX97fakz483Be8M83zeOOI9B+JhbscwNxO4TH
4NSVRPRfa81MJ/nEMR7q+Wep6v+8914Vrk/wYs5//W2SuzkmbHfzi8Xo3+RtYjTUgX1ee/MyxkB/
qslC9B439uDZhjxdh2rLVi+Z1z68jUDzQwP47GAAmIGJUUyWi6Bc4rjHLdElH+YvGwnur8igi+Ja
7IvCx6lUC9VzIRkiFN31QXkMCuDKK9v27VeZWCFQOWiB2vJ8fuF1NQcZrQn1jguZvdH1QJ/RM3Hm
y3C3iYp9gFzBWDqPVEtOpyUfSHmcJX0iyUOU/is93BLpgNc1YKi05AebAKCXG2zHwZJAyJ0HXJms
N8DGDcECBZWwfNvfMnj0G6bL7RksW2Z+aLKGvSSoHtvcphgh10LtdCkxpH2bpGtA9qANDNnWFL8r
Bm6FBo7EN8HwRFx9Pgi7LppJdv3WcMepSADFT9Bbu9AFQXcSsqqSFchaYVbu4XjNGixp5cX2ginh
ZxaEUkaTWl4hgn20xMPgnrwlvjsQwbIXTVZlCiT0UzDULVnJEfTSJNhTJNRAenoWqgFzIIp9eNrk
FuvjNPw/nCqpo/Rl4p3eH5coGHRKlG1asms527w5tW6AR9unlqqsJCIaXBwqdz2hwgHC7wR4l2V8
2S5+s9f14hD48mkFd+7YbH1uib1dtqqqWaiOec4OMF4SJbeBbqDhGdd0nUtNdnO9lzVvvlCrBfZn
01koxkAPzA2WKNPwOt6UM1x0NMlijrbgz7eNKg3D2NaOZf+l85dsNdPYVyBITkehafXc+sO2tIGE
3LYoJ+QHBx7DwHgGSmafTUPC+uEEy+x48/hUNuzIxdVzJ/Gsc9NRaNl+TP1VhCcOoWs3FsWCiCWG
IzatsjVCUTAq9EMhX/JTJj4z+MzC8762LE4r+d4if8hHF9hen9WVWSElCjMCwghuGSlXLW5S2CTY
1xSFMM7ntzzXkRAeAbpi35V0ZSRYZdi0bgl+cZkL2C3DmyCWPtj+vUirkvd558rKhHV6rtJMZ7DA
sooVMhaINCR2BimBFL9MYB8OZTUdFvsADIV0dkfTV9Z+eo2HvNyABSUqJzlZ7yJHk/2BPsKzByX7
QOTCpHakFHt39ix1lwzvpUd6MREOfqHx1Oku9zLHh6w1lH7S4wWynKqCQfCnKB/tPWYiiD3tXo4S
3fp9mJPnl/MD7GusYFKjczaGcjF20YT5p1rkp90IQhORj0lx6YQx3O3gxqRISWPO9PaLIRI7JPeH
HN5XFLwL3X8DpelVlm9FJ9cYCJVbBl8oJCQysNrYBD9FbIcHhwDkb3HInxVIbk0h1+rl9ZXkdIVi
2UFEUHzSxpy8Wn1lYIHk9OlzlqO61GugrNPkCH0X1lh8qfMBMD1JHMIc2Tk/MfeGp2mXX+QUZhey
jejueAKwC1YSj1faSUtiw3RAF5nH5xT653JTSIbhFqXMoFD0BRZvqs+i4OJXFosFbTaAcnsj/Zlb
JopoLJ1rapFNX1ZGqZQcwmpTdmZajI+W0zqQHlWzGNVh/JCZ6FqcVr6hZMTK1FmgyVG+qW5nCPkB
KJI4J/DCeNK23wQbGGPNa/ssm/jTS//sw0aDR2Bk8yqxwibllW9VlJ3m527zpyOmaa1d7kwIcEse
xvTAXf9au0LIPs3IonWR5CU+BUdl4Mu4GerWoJtWuiNeXR9CNpuKnvcNsijbKGxmRBdKJfDcSiwH
iJ82ZMgButfj/M+vR93wefihQDwnRYzNrzVk2JT1oHeixvRg7wvpyFxCfgOpdySPTWsO3u25Dgzn
H+ie6NuXwU3VmN/qlRnbH1WXIjKejXZJtAtOM5gjSAbwP77sJXYIS7BSFJrbUn9qbpeLUqUfUmMZ
6pVlGTFfshwGMLbqcDIC9rktPHgEjNWnbv4a1T9xmR2MTHR0fMtI7yUvuyHzEVyV8RLZt3GoEu5n
mZen0WFjN41wr2XY7x0B3jRrJGMljaRFBgvTQ6uSODYdibLgNPXe9NitmPFt2Fa1v890FttgYgUG
54xSyBb+QQpsXr6AV7lM9ZaU79Q3AxYwZT5t3qyzS+ExgHKDEcsmG7V1OuPD3xIKb9VTU7mPUt0p
jhXGW3ljhAvkYebruYqHpQ0dIoZb8p7GOrSzUP5c/GHq+rfNygEh3LW3qhA7s+B8zi47hz1bWZK8
ETMPwRYZRDfWiiD7mgohaVRFgYTc0R7ndokRTAuJTvpGYVxHT953F6uUQbJoHN8a/EsuJKOZONYJ
A3jVoljpa6sKV9uPiXpJZvdep6fn5kRr6k3YJGGMT//EpfPdlDLg3FZcLN1IiE5Klla8RDvjESlQ
qqqS9hCt1ULPMSfUle6EFRem1xNHGBbnBwHXmopok90KcUtKCH9kIxtIC/oHr9PL5lKU5MOEnXhH
82f0Tn7O1k6DowvM1RZemY2LoSctXRKFfSz8rG3N5QbAyNBu1vmoOEVcrdnTTe9jCATljJaAfs8R
OOnCHbGjuQnI0Wk/gDbXBv/Dgpchewxty3Uqw1Mn083QOjc4gCWb3YGEqj7j0dk1AkIm4etirKKi
y7X1WFc1U23XMJVyVPq8eunXNiUqFBJsNPq+do/E2unNjlbp+o3KaVRpBpUWa1EMAaASqJT67jzE
dV6WHi4zg8iJawhhk1laiH65RZTCGSL5cw6gXxlAImFUZ1bT813bYlG/30gnjtunrK8w21t7+9Xz
yHuuBI3V2m390RqA6+Tra0IW4L8QZ3Y/LZlbu6109QrAuRqob+/B9dDcpqDGKYbrhrIYwJO1/dB4
WYHttUvbOlHISHaaMzwMiDbNFtBGd+34+3O8Vl76CXmkgC7CGtU/7fSCjBvIRlO2ZbblXibMkuWt
fKOjMrQ9FOU7LUoat9PY9zXSSG6edmSJYlD4wC6V3OozEDJu3yldRHUf/l936mU6+xod+DMaeVQL
EGZro6CTcPTM8GN8RSG8OVcCwpdL7xna/YU5naJJzdreQJ+jIl5nMyx5epR8GxLxodbCfl1h+FTb
Qyl+onEAnVH5PStLgcY+YNmwdgBsdv/FLuCJEuXtUJuL87j+vOgofEEv2k1mxc/uGtTBKsQ/tDHM
aD1NrKom3xrSNsXDFPG7eHFfstVYsjsbZu9CW9XKwO5DPErSsBEtvLz/dDqoyDIiUI1t2Cjr7y0g
uJa7SAWYBHHhiNDApS/fC0rveCRwqr9UKvEYlcfvoXEC3i+HNTK8Af8sKb5BMmxRdPmDxyMbF1TB
5wLvjXA9QYDBpjQIZOAMxlorWu9ZH/7vIrxX1DUBGPGr88TsWzpq9tk1LStWRv3NJopus/45UWjT
jA+gg3Ez2PEp+gxerbsoUwFjN06ahAjOU902wLecAkBlV/lqSnldMzOwW+iqwQ3noVV46dfoOlrh
VuOdc59Qw76q1OwvP2SODS/6J1GD6B//tb2F3wpl7WhlPkWEIFJa1rRg8eL6iI0pCs0S4LAGIOIT
YUCb5n7V+71eH64bZoKN5AKLxeohY4/n0YXVPlr8/DyjKd+QTwHJFiFaTM4bbc6TRn9bceFUSyav
7fGpieI45EfmYNBN58ZQxrgvDUNWuFQqc7gjUjcaMeTrRfaMwZJY3PKPC7mbhhY5x103jy3TFrVF
tASUiW6zq5bBlAtcMGfLCCn34Do2z4hNLou24SQrBimltXvFB34zJw2NwKCrxHt0BtdLOjkVq1YB
RZ/lyVwXFzRFyJ0OwTlQM+/vgWjcz4BV2+heGST44+QD5LbX/unYJrwhrCRG4U2IqMVdLfyV2jC1
QuqjxNUblipodkgy9UIT6K+Z9mbdOjNb4o6++b3EcKM0kOS/bujXnFAcsGhzMsjWd44RSYABqxlO
awXLFPFb1ocxmU26XQUVeczkSn9LvRwJJwu55cHzQu3N3/Lb3LnPIjv0Ha5p5ogMHLW/JWiK9Gf3
38iiJ05XWD41VxJMIWWV/OhiGMfBNWNyx+cyHi1yxxgPMDpThJq77V1TIHddXvXxe4uduMtTfElU
9SnfD6Vf6jvUo8R9bhG+AA/q1dN7od00LocM6kIj/IuvbGBXB2LMjY0q/vyLfeIj6950smPdRl+P
W/JudhZGHTBFbseyGtIHGxr8KX11OE7ZFBOGRMf3ETNY3kClgywxVPtHPmtdfbsN2BsaDLtpxok0
1/t/59h0WBjb8/U3P9lVFti1Q60Gp8s8NctBwvs4t35kdPhwsVIjTUGyP482ejaLkMsfmwKafJ5x
E+d/jcmYkcx0v/YrMbRFOiSXS5vn33A2joOqeBxuabpQqcF2L/81WEirfdYYREAC3M/kZ+PonnXI
Zo2QTWAJRx+vNDABTvQAzngcpeW6KVES600dQXIBXzqB1+evPquNKiZRG0lhNHHtbzpdMuigEAH6
2L/iuENfTKb/FGlQXc4IDZUhIXyigSiGxr6BzDvUGCeZ4e+EbqwIke9u9jGKSHZRHF29mLT6uHtC
OdgrTXwWqaZCQpR+eVHqAOuzKrRZ2UsSV9iH0Xw/MIwGCelvJw63a1tmIjlye57bch6UxVO/gXYJ
febKbpWqh0KYVcSIXpGQ7wVGrxIQSpLBBhjNn4OQ0Eyu99jJhvdFNZAGEAcTqnFSycTS5ubIHlbY
Fi1SKy3B9Se8Q0hPzAOK2XwlxZgtj64sC5okszhCjyOFnGBQ3gqQL4GeI5Jspa2BQJ8eAsh8EZFo
gzXmEzqNNnEex4DSDNperWJZJ67EW5ehOoNjLqLsIE9SI6G1xOK0o0Ht/4ZAvqJ7jzHK24wfNGkM
e32mVTgpA0CabSgqFFUXAPwZLrX+cl91ADfECEqpihywNoQkXfZztMdV0htHPobTEOpnOV1yn9WE
dcZOVwDKJ9nRVEMZ+2zDzYM0KlKUrRspg0YqNcVDWHFOYaW9ARRt4JttETYczuIt5HeHoIluCzhU
cWDFqpEkurLbl2F9QDP78oSmxjHZlNgN8ZXyJ9GE68+DycXFvFokWoKUyjlpBtKx0zji6zs0DBPj
Sf+vGFQ8CuSRrGYJsvQA4KOZvTLvUAuKUFbnwUsGR1Rr9SU7N0aACwYkpn7EQAM2hEu5C1tvgi6A
3edNdrZssQx+sH1NRcHGUSh5Chp1uGi0Rp/ctjGqzmXPS1Fr+bGSHGC2sXNWpG0djLpC0lJGUWv1
tiYq4uj8RhXJD6NR6tcEyeS0P/3jYhwL8N8PpDlxQT2FaPvY43lulrW5N/vE5J9JyhOBXWQkZpkM
OsZDmR2zcbmgfnirbdPmIKZe00ktRvPu51YVOokKESkHM0byIR6eR+AxsTSmFjRYgRGX89KGaYcd
WLVF96wrct7nyDqZX9R6rOfTl3eyEwZ51NlMUkrYvQ+u0toAypl3B+7bqzAqVBhqn2jQVWkuLF4P
CVfX7yQSILbE3VkkIDguyKiyuio4wzUZFz8dJRUiI9QIeLjoU/MAyacWfRbJZdrTXMWuu+Hw/yTH
WI2VFxxFW6j5s6RTr9mr4uqR/YsiQfhHJ+RqCYkk0TIuWlRkqOqvpcvQ2MEnVwhXPlydx3BLXfzu
2Pv4yddYwa9/Fek0KJh6qFQsaAbfBDytKR2qJ/p0KgU4HEPDI0SY9aZpjiCGvEbIaxdAR9wsv3RZ
iWd9jy4tm+61Wo3HpMzNYqC+EZ/fZbDn/AmpEyLJ3354l7C72VkeIslu1X69xSjhsTme+6zLg6T7
QXlLAe8fjX5XToFE9aBTIh9F7EpwWL9xuI5fpXTFbHtE8b7tX89L3bZIITSahgXlH7WFg/UmeNez
zpwc21L4Qw5KAH7+6KF5+C1Vz36DRJ7aRAmW9MWRwA9GHXeCwEsRXODlWC/ZPWd3ALViG5qlJLnz
ywZVhgHu3kGSMOxSS+Qgg6YexR+KIO+DL5sTlrOJ6pg90kbj+9QEd1llWPddPZ6cNWev+85U7crO
TeNutBncLJ7t5oBOLoeF2JVV4QoQ1PsOXysUG8Qc3i3pbT6yzB2XKxctaD5ta3F1fOd11mSKcTBR
nhsi9fPqcLyZTMFqiZq7Ia7OPuG5g9qt63Knq0d2VqWJbRuG10CX21cTquv4XWWb1dC2e9a4trjr
qWCDWwkLXlVJefcIlKCDdn5iqgVGvpGBZTGJdYhLiN5sgH9s5pMngPVcA+IvX2BrYuSaby05m+Rs
gwHBQqo2hEE0iSOqdqFChwxOEvfVTk6qSzZtc3La2SMFWfLOVoMbhO/PeICBkJMsbs0nmpn+Xxgm
Nvm4f2oiUDT2J1urFQgoBRzebbvefYdB2sLA+sjyxuahuIxIsnRbOMz7VuDmG/nMyLEMKbWX++pc
oUf71FZlxhlbBGRbv18Z6XoIA74fRcATlDsx4cKGcy2oz5hac6DdlFHwD694uWUdux7QxxBlbvlb
rWwTZ2TmVQ2qVW5UtLFDr6rKpLmE7E0DReQVMtvGha7zaAMsGuFN+Ko3fKFwhtv49wGPEn6KUHPD
eSC6SWpHhFZpy6CZybg41fdkcOozd27E9ZgfrvLuk71+Dh8+4xJpoikPORmNme72NFAfdrZbQbn8
24LXqycbwdTND43x8Bdni1sHtUxZpDoy8pN5hLKlcVSbfq7DoLfF1r2rtxJ0zxIIo3HS+WKufYL9
z5C7kdOFko8DPTcMp52o2nHnYbi/FYR//TrWU7tz96Dc4dKgAdy295i0YUpFi72xF77Bh8d8uZu1
ZoKukvuX78y10dXBCIaGwMU/3KnZbgEYeYosJaeW2brcDyl74QWRFz9Wh4MuQWdKfTqPTwIoV21y
v5RROkwNxJXhx+9wjDqXOgjfhIgFI/Q/6dz2CH2moQ8vq4VbiWdZaCee6ozyR+18qeU/B1IxbKDd
ONRoy587P6ntzpetnJyR+zb6RFVRR0rRuDQyqc0X+Q3kNbcDyXAaiCtWNAM4NZZw8MiUv0Sa7jwi
pIcDKSQzhyxVzx++M0l4DZQ2VfK6T2nIFZ7oW2SajwIfXF9FoYt0de4XSKw0qIHKPlU/xBdq9NUI
OU461dkX3KA0UxCoKDJ+IhKJ5BFEbdSZk7iNqqQk2BvDCcrHc8jvhUGETnTtIxqHXa0qFhFZYGFG
jy9GKh0pOV4rTvwpQFrajQ89yyAUJyO8+P3UX9D7mVyGKOaNS0d1u7ct9+gRsAdZa/WGqskKXUcE
WTtc3ISEEe4mwRxMYbLAFIil36xarPDfv3Kl3ZXpeZBefgR+3kKQSTLGC0rjgEgOjTMpTiyQUd3z
uThFa91BvPmqjjA6ZsxsdLIT4gBRNEY/F9pU/ps+drNZxgYIxa8IMQPUk52FGh6DfXarJIrOlLD9
jwBy/2+AE5WwyaTTK9UgAz/mhkDNffgVMqz62bE1pEvsKucdo/w8OglghVRHgbJvNyeiU6YcQoiH
NeWGmoQGO6awQRL6cFjT3O2eJYR3UJ4Z+jYeufWkCpUnyhge2MF2UGpSkWZNukCZIb9Dqbm62pXH
xFIPFzobgo4qfUT8/7Q06nojb1ZhL6EgzgdWQRvDJSfpP5JlwV/USpA6PsKlFkFBhayQBAm6jzNh
2beuniH6YYfE8KieHYmyhhl07vffV8GPH4rGG8iiDDo9bmpa6itMlWCt03nRN91GrX6IHtCT+ACJ
xQqkVZgnatrhCYfJtmmIkOmZQfkZvmfXJ/6nr76wb5YASDOsMJUULPLG7b1TdCdEXpkRKVJP2gx9
uPOCUwpq8hn0F27YKAJwCuPH8XDQBcIvysSyFr+IUE/TKGrlvslfVZxjRYJKl60iHdnTW7ZXhyeM
y0B1r5wOTs5PdVX7KM0HMoEU6jMoee5d6SF/YMCY7zRJpJANv/Jd7LIRw/qIHyQ7gtHZfiWvvAFw
imSsJ7ivqMO3mQ3/DfMHPqDGBtC60jD9LdNJ2EXyV9XuAAgtcaMaEGZPhKCBVKlpIi3q5QmQgNkz
6i5ZAcObvgc+gaE3fmwgEHDjMbbleYlRv9IBikyOJ6ISoTBTbTe3T5EhvBeYJYodD4tJZxvIeqrd
37jr/Dc4ZXwar3UzwL2pdbQM7Gk0y2+ElaCZdJr139GExTZ8yKNdjiS+NQ1d+UoI1qOejIALxWga
lvMt7XYbUQJlwTvaJd/2KIKRRSo2yW8nkRsb6JUhHog2Un00sKLeqUTt3kHFV8OcucwOlXT0EW9A
osplin6BSdAqiYvBWO5fW1penfdAY32SwyoZqYuZvQdOE4cO8sV/XrnDiNvXQYxSsai3xtX+9LKt
+kKbM3ci4OnJOKahP+M+h57r2ZuEia9v+QQjQm9izlHEr+uhfsUphJy/WeHeZrxl89VLJP2Qk0gi
Ef+mNtJqGSKShNxwpN7ABdSw6ciRuEvlNeLw28F1Sqdi5ODlC/GD6cDCMFrgn5WYXYNaXJsYNP5m
rO1GhFOv2NgOBiCbf/arTnJzE+gRfFckzyJPf9+q+AU8YrXlvSZHrm8Vof8HmfMeRr2jjwgCzM9p
GQ8l0HoiO7V+i8/1hloyKQCAoUHgc+nFfZbfHwhwLjkoqqiOoDPe3iHk0SnBeAvQxGdplVWbM4Uw
quOk06CAQ8/g8fxNnYU7KBRu0vLCf2Pp7z2V6Toh8K/OiRkVuJ9F6Rxf4YjixW0wFPEpC0/yRPoA
uvyHEGp88nlZsNlIDWnaGFWPtxLrnha3JXMi/IBWQQyhqdYwErlvGfbsdvrBDweu4GHB5S6s9OG1
Y4KwX0eDTtSOdWThfZ/bgZUDLaYBabUkh91po09KG+/dkDx5mZ6yVmy3va2DYT+FSzKRR3VLXtsB
hXdaDzuANAmJGMseoB2WnOxngQvHpIQqP4tSGPUWDxVI4EJpl7PMroWv/o4uAuH1dJq5EcBY2G1U
YbY1r1YZc1uDTsmr0RyHXv2W10t4w59utYGG/rXMAXHmrd6irqVlP7eSL8wBK26BtbkM9/nKOn56
W0FF9WFmZH1W/3hkPFPSt4BMs8XNDTlagQDY6XSIXmVmuD39j94gCkFugnTisYXT32PCn3gruSX8
mO2Cvpf0n4CadplKD4n6XBkAyAokoiJjtUPQYlEgz98lEfgtUIlMdfJuZRiTi1orkBlJJtWHdZSV
YGKxk5joKhH1w1s/ivLXl4OXOXw3KD3rly8ZNfuGDhKXzv2x4rXquXsIFeo69dTTcHpqnRHXTfd1
3lnmZ2vE017Q5CXfjuLD1fd/aLXAoFSPhwP6IcpuePIe/hBnx4hnPqZamHsF1tfVYNg+htlT8RMz
jeJujWhUa4t8H933sZxExypDC9NptUNYnyfdR//ySPwasAXV2tZTgcZr8ERPM32yVINtXwzZkoLA
zP2c18cAaP2oD/Se3vVhcKL4ChgKfJAJWjFG1kui/5p93ZaitZok7/s76gEelSrSxfzmhoTfYgiw
YDhjvs4gE9zQ/0KaoB3eL85JX7GuKEF8CN2S8QkxNVBTLIBJeke3EW2mO+tGy9EUW3otFoQemTgt
vgNhQI6z/LN/8a/MOk2S2Sq0iH28L3viXpkUrRrXPq3r5NG8lYm4TvbFGStMUYbYI8IZjvMWzZeW
FXCa2ASbJbxy9eJOheJwnjc1DJfvJYj4GZXMBh9cHkaTIlQx73n1Vkt5OYRCGu7dSWltNvsEPYIK
pHv0gUS5XH0VJbt2luq6Iomp936TVhMZK6/RwcwW49y1YXJ/0iIHdoj9G1vB6KK81sq+rgITJZdf
Kgk8RTyf+pd1ivn4KyZLm+Ry8MSo3WP5/SjR954rLEXDy8UUBQY+Ne4YOy0dy6QkSOFjP3AljEiK
jG05O/xrmM8vhvBzTtzmP8PuEat4DEKR4oGAyKl7SCchYv+d85J8ojncBsiwQcbRdfiqO2JuCLHI
zVfE1v+/HJo6+B/C311zfKmQWLHkjSuuEns04Aufl6QpddtwpTBnwDxj5l+CEt+Do6F65RRNHwKo
EvTp9FueXZ03wgBVnqDyyD5+fjtS9PHP20YQsCZn9FOcVaygGCdC/gtQ9ZZWoAnWVhjZPELt51ii
YSzMNZ5RZh0DKhXlCqnstINW9U4jZHOGvIDK+B19HJDxNFu9J04aI5Nw5ifutzbpFyhwYBy+m/6s
KbgHtbng1MwicyQfyeuSZoXU8bZhh1hx4pnNMrFkfL80yBnHjpYIrlAPSrni3gEpUpiVKkzj5Hzg
O5ukkol6bKThbGyk0e7nQszbTDaI/pJI5p/Ut6zj+pdItlGSnBCrdgyu9zTWKn6GFvuauuPsOlbc
q87ZERCCsjbWcgoNJK5uw4RImNahcBny0SBCL3e7Vv9Mr/apKyifeSKC9/t56Mt852/huj92j9Q9
MtCyIHUVA1b51C+VZe5CkkcVS+RmJLxwMZmAP2AFnOf2twQzjbsOvLgqy3OkJRTH5T6oZ3cTOg/u
4Z8NT4wrMzHBnyYTTfEOee0NI9VufuOw/DbDABEtYnK8WgYXCiuhZlcnaFxAM91a0rVyFRSnIohz
Qugsjq6iF04j7Q+IYTJo1yhxjmy5vIPqj5Oe+qFMUdrcsDocPUPAiRHUZDsTd169v/mGjoKomj6o
48kwetcCSo9t08GlDw2sFkeolpYZrV3+VrGZvBDnxEP2pH4dgNrTAgoP9JgxxjsjuiIB6fhZjqV4
n1NVPnn4lMT0/qyXc6fOUUk+cPNg4hkmjG/kofGHzpZlO+/KG4Qc3W5hDlqQT1J36L2DD534MSXA
yd+9ODPF+23p/6J0hxPTdEGG1z4gVKA+a11bA/oC+oOflg6HsF6WyHgXlFLyfi0v+gXpuK5ZhBGE
YmUN42MYJ9cByoTiPZL+EdaiHFuTZ6PlZpuBjeZrtraj42RkNy2ZXTE5x2znaxOTO7wyV78+u5oW
fUrZDMA8WivRtfjwL3merNdNNdHT1otbBg00Z79rO9QUeHIIvLHGDFemuQJpGOZPK7ZAOivYcD1F
wv5IZ6bJ7vKzBDYYLWOtlK0bel5BJN2fzlNm90VbgO87bBDlKzvMHQ11oz92jLKh1DxBp61HwhSx
u2Chp5Cy1f7SbFFgBBNqfekUfYiJ3MHmS2Ud4aBGi0DqSHAAWuAw3IEWHoIqr0C7sH1UKjLlztVs
+T7nB0vOvz/VqqSMdpsQ+hhiST862/Mr/A6Hua3KVxSO/HciwOB9opBZn7fvMo5vxzyU5d8l5CvZ
TN6pvYIheie98UeQqznrAGUy1G7ofwH5hkQY1ZOZhqOwXgKGyX6MKcNNbhlWZ39lfonB3sjXi+PT
ckWtfaXcV2QuJZlJsjoPS1OrK+mo+pRuyqTJBI031d0tBjdkJbm1zVOdKMDjXVZJpW8GBco2z6Rn
AW6VAkgWo8xv83mbdm6T5uK1Ao/RfsdSPqNcit/E3TZ6irWINcHPDKuFIblsNK53UAbJOhVn9y63
ZuXUVeC1Kk7SDPwmUO4MbSF2fj3zhz58AU3/rqCKlJE51e/UymcMOoFlCHlkoekS8At6lZq805cu
ZYVtc9RWo0s9JpH0me2XviULdCPkQEpEZ9oHIxp95ylXY0MeLrBdEdID2nwFoD7bHFiOGy2DIi5H
RXyPELD4rAyh43IB0NgIk9rQl4NIuWMi5gGlI+sXo2Whyn+HOzbInatGc2+G1HnqyWyFTBm/ETsw
vb0mZcHomzhETFVNE674bcvd8PwbaOiMTLbNHvsvRT+d+0NsQe2hYW3+EJHC1wI4lW8dbWzRxn5T
bf46d1rQf2OICCFrx5t4+OU39RNMKYBlSBdKRjJ9ODsklL5q8TvqbPueDhTvrZ4DVb0OcgEb6nOk
PfOdjU0FAfNubq1Pes1MtH2ySm+WSLiVWX0/PWo4/vUYn16PIcx7QvQsvR+/Y+2z/Id6TDjbzp0n
myZXX17CdigACNPgBmLeRxFBApBGz3xWDuFqRh7De8weNbY6XFKGvjyA6ybz05WAMfhbTIUTULs9
CpbzYjDT2H40fQCeIcM9T7nQ+xLz0olQW/lmBI4gpfxqzb28eKHHG6FkM56Ln1+7fRTpemGLD7ai
6KSKhl57Q7CNj4zSJnP1AEoCCvcgJDUFKwXmYOhsyqoNHThIwxnZVWhNMR6OmvGxXpWI5JQBezw/
7Il+FG2fG9opXdzK268Wtd1fOD/IuWTEjpiLXvYE1WvrkVqEo/8TIiMC23E5K0GC71feT6Y7NKBM
4gF9oLraKRvDNURRNeh+Q3Qz/UMYIpSDrea/9DqSBMjlDhR++JmCA32BiVcoSTeWuSKAlMYEL8s6
Q51zLwXPnV9hqrqWB/N1OlB7l4+oGEM+Wp5hqMlTwTfIO/TxGqww4Y0m13ClB6o9JlHWCLidCkBa
9nPEbOe0ejVPHmMWRY572pGm1o3yU+ydZ4Itv74VDX4XnYEy69Cc2Toam5Ka46Bo9nZ6Jf3zLuch
EI1MrRTk5wsNTIqBKGMFgqkxvz9XBistJxeQzhbzjYaZACBaCNaSqY0brjCrs9ULGi5Lwnsk1QlI
jtzHx0CSbGK2qfcictzNXbN3nU1t6X/7ynB2J18mpunQDh8InVNIU/nUnCKcM6Nq2w+Zf3JhYoS8
7ltEZRtYz18+IA2d8gZXeFg+YZdkeWAfdrDi5Dmfpqccx2IHHdICWYzz7v2I4FsNQc8hVYfeH7Iv
BxhQMWr7kUND8iAZOTrOcpUlrH8dnrj54JsLoFPrCb/SYJCCth+dATBKL/W2fws78xgEeFB4NeEf
IOZ2MD4/KdXN73xNp0M17fXxyMc9I81xaH0uK8TQTAdKmK2kH0La6ALOrzKPFQNIAA8Q77ZuVFkJ
bHFzgw693/tuzj39OhZMokKwe27wzNx++liFS27Mk+bMgW9OI7qESwz1cHEWQ2QaaKQvN8HX4cMf
APFOgFWiDomXE86V7iliUSTmr/ILRO986m2eZk9doK0yZP5yZO7i8J7mabzkFfw81qgsajkwArEo
/yUzALQTLb+JL16fzUX3Gww54amkll/XqivFdzr9mNd7q3+q1A72eKcQGphW0vbogKaf08zjMtjw
nHjNeyt7j/YlR83A8RKXuIui86YjQSITmtgHYKtr8ESe1yD+TSeMRcGuRxcZDog5wTpmsJnt+Pv5
YVPeGn3PRsYq0RxziXjguMIIHlQcyl8f4vZ4KQ1Wrr0MfP8ZmOfTKPkTBea+ZYOtPrbQhhd1NNeR
XVW+JRAjulrgzRTLlYNEg2odrukk44DKYTgWJZV/fW93fdmksTXTmVLowAwo281OmhCEI30gt4Vj
jGyhEyNUB9h50Uy53Uj7gGOiADcEa5NYVlVfZ0pVRLkN0ukSK+VaOc+CphUdUJmEyTie2D16yk/l
IMwy2ejf3Dqin1o2DgSIeEa+17cPfDg5t2Pert2Wp/uRSnY9OAEOTKMQ0K88UkLOYmk7SaScxLKe
6vXJo41Zr9yRwKCFhqVXxQdUZ9PR4/d7HXZHYPL13S6mvt48Wy9j6JSzCxto3uKrVwOvq+P24IvD
ndesOC6QEX0uXRGe+IiamG6McFAYyKbHsQBWCIyADe7wW8wLd+9E/nJgvZkjNER54GbY4eyPbnQf
mqs8IWKfHIkMZMBXS1n4TeT4DNdWOdhnB0V1mdklSedjChUvkpyGwfGn8czWlOQ3tDww3eBVjVfK
SPB1hDFn8Kjga7eIaIJxF+5p151O9XVbu940fIrBs5LVLCKgVfqZsAv2kb2D7lO70wUx4a9vIkWZ
YWwn5TvGZ1B56bsxBaxXvHkVvS1c0v2ZjYgFRf/bZpcVpCfUuNRDpuSWcBsnGYSGh50SxMvOknp/
7F2EL8cbP7w5ktvtDtDhFIMtlQ+mQ5BIC7/1Z2AjUeD6QF8yXKdfM+Tr9suEDp27KyfLrvY/Bdys
+jDdNdoj75aT5GHxcvCkrtrQudAHQ+V5OfIwp6ZSDr7mqRac4ekZm6OXfwjGJBvCz1dT8Y0QWL75
3DLkr3/6DKmcZ4yh/ZL0Xtha67t8PS/0RtADDqgD7eYhhwYLhnidOiVyJT6QADc+W8Lnt/JbKl5M
hl9K5ekHU0sRsXVs42dG4ZC4QnXHPV8pSt9+TP97FLzUGocBJa452eE80kgu09POEu1fmtSYV0TU
VQJo9cdq65AhNUzZ0mfqwYvMb+He11NAM7rvH+8sO4dEOeDJSAeoeqKMIvM3xIpBUSJyURBqlWRi
cyFJfnpDUMPkgkRwQesJrFYe8QVTXWDTFbHR6qdGQvdbAaJVkQMgyK1XB77r4bmGwG0mkOd3/H9C
Djcx6LYsxQ81MPDDYGZnchWoinmftluTozly6Gk9NT21Hx0zGMHD8RdPbhCVQKKJIShqtk5AMz2V
vSGPLXEeRGIRQLCNjQhg/trmTpNIhbgXUVJGQvWCwOJDgRc7szhdWPdzNveMmU6Z3rPlmqnDQKYO
Iy/zCydDVAkXRaZE2/+W8ob/YxMVOTVunyAjmjBQxKzpv0mXvm8AoCU9IPZFgQBAwCiOG/JLnOSQ
KfMNykbNtV5cSDctMEK17T8Uav1ElxQ5HYEo/qitP/kq6QpkcRVaRgv/xe08/w+MmPuWOeIRjboQ
MVaX/6iGOuqVpUtctvKdF8dKkeeZcSuwyDhGfsLRnicNkpUEd4K0XG/QvXbdCeBimuJ35/+P7/GA
8bGyE77J2nTU/UpSfhuZd/CcGpKgsL9Q0stMaIQwAJ9QbDNe6lSLv5DVpSKPSEocwR1NsBjIG/jW
34kkmzM5bhFI+u3Yfw+qYDAaehITa+R94qcTwDYyFyqnUsOa8xRg5wChLIwqIYvbfPeBVfBgNPjK
uEG7tJ+EmJbfLwYT3d1/O+M0/me1C+/AWl1weyo23GUxTglaKIfD/fdMrP2VKGcrP+/tkbI6qHCP
2tjdQ9JUJwc0XfBF2kwcASLC3fdE3R67ofUp+/cm4P0WXxmVC3y9urBAgXBbQSLatkDgoeqLAkpU
BdhnLfbctwNnbIgZEVmPoZjRGFvE0vV9p3iR68ZcJQG0vLWRTB5kBTfITeKH0+NO8oXEsvH7p1RY
3zaTM1GgmQK3c2U+m6IOfBGCAoK/64m7Jnq918lxr9fz60bXOZxSaoSFXSTh3tIMySU1vxlV/At7
M7YvXrUBsPWjMydBihNlARXUfLbHYwPWo38a0823Q9cDsG9tILEl5QmsktEtARys2UBJFtgnAOht
O9lnA+3dCuiflSW7wOHLDmgCxkpsBOktazsJg/2Rf/mBPOXWE/2tzoiEqs+m4shKSNkz31KHH6LR
BJVG47ZGy1w+0GdMhjmkCLX4bJ/4Nvgf4FC9FJFB8QQueNA2NQggYPwT2RLkb6eVD6jdVRMGmoeu
HlwyqBapdfvWX++gRn/6aesiNIzAR4S8YLPd1Rlnv5nMFD6B34Qdb+feEyx4AnKNhFetJEEJfFyA
kGYx2pl+nxX8vdGLF7xA9+NyFKMoBUYbY6Cl1US9J2xpJWzyFuafkp1+RnoIJkv126ymEZCmloYJ
35+GFlukjV7fDFYK4aNqRIwDUImAN+FdTrUb0MFpIhCwKwDDxK6ceKAScJuXJvLKoSI3YSUsda2A
DCrcd3H5ZLB42PbPua8lSNpQm7pZpkA/odc+V9ENcolmVSJq0jxeaRcF8xykwpW/jKoxAtxK28cM
qcdLymAsXaVhYWSltRGDJRlH5u7u/yM/fMYXxa9hqyl0EAS8FaunoBqkyXTxXS6hyjQV9fRluJZT
6QH7Usx9qKxyirPdgJMQSxtKYTasLI1vd1nGTrYHs7bBeViqJcRlt+87BpMPl1NDuhJAIamRswo2
qqo7ujBqiZokcsjHyHUVY4IHSZGsrKcj6fj131iQ/h3xK53GeCXWAcTETwqA44hmYyX6g5mJ6q3K
J3XKaupZYukp8KuXLAEjUcbwX4Q4hQMtvBUkD+b7zGSpwuHz6mTBqh6wDBc7c+3WPxguHr+QO0GU
EDkpeDnFo8WXAXFTh231ez/5NFqwRVxhRlVm/u4axxLjeydvunXYg9rrXFt7XlcqPQ53jbxk7orX
sFpJeyWu/2eKRtIXOFkZ7O0VkixaPlIsSwoIxIY7lqdZMutqsWN1yPo0fo9QPDgvG6g3Mu/bU3zw
XpkAq+q5U2wQWAlh+aNQ4/vZvd5VpDictVOUKEOkoY2CRNHFEvijlvkEFB+EfeCIaUHFgVL2Lfni
Q7oRsOXPpAUTcT53fy/XJVT66HfV+Cne5Tl6KpK8tNuTZi4qMVM86KKlJHIFVvzL8kcOiCbufeaL
RZqKsJs/7I5IRvZxQGHfk8FbOqlR9ZBXpSOtgzJ9Yf1fTcy0yr64zPbS11T0XE1e3e5mOkhz4BQJ
pWKWIduycXD43wVKmqRCPP4KX+ZAl9gTYZAhstf/48aDv2sS3X0Zl37zJXclxgOdPdkm5P1eIbkX
wqEL6LNjoIg9MXG/JPjT4ZzxwLA6TbZC/EYahK+3CBep8AovkLW9wYb1az8uk8OYXv6B3SxuXd3m
vMOQxvWAiG6nYr1HjmS4YoXqwSzgUvN8pIcpvx31IbnusU4Ks5PRJDWE9Kufp6XgBMA5Rz7dIiie
ygfqHVoqCvq9XR24zWMDBpQdfgxLgP4DP98U3yafi1z82Tr3+Zb13MKcH9R2YY4D5XnDAvu0LdGj
wQf4EkSn9yvfR5wNBYOmNb3UE1joP3c5zU6n8wSBXS2pXKswPU3+Zh/4xzmlJVVVFM6EW0Usad/q
k03zeCheRmgBQ0Vk7B3w2CO4pqll1C4se9EsINrmfncb0yyTRXzi75gCgdMLe4TFY1wApO8BZoZK
eUtexB8uYoFYosz6aAxDC2pvDm90A8ZEf8Cho++c0xrMAIlJ6BI/4Tu5jQZ4L9LsVAbCqc3GovSO
VwK/l9v64zATsEp8QN3hbfQmzf9KNTMjqzr5uQNCx3er4uXYdUIVbwYXvOLONskEH5ot/ABBvg00
QDUNahUmalzwEJ4NvnXeXRvCw6IbTrWNWBifJIKBEkNU4HGnYKMWg1jtrllBmx4R1cZo2P7C4iAu
o/WMquyUzz+wjEGpw2MPCvsaO/5O9V6uBq/qgYWnOjHhwGkwz4VnZgfFVAXDsipACGCsxgvW/Xoo
bAKhDKiajt8VPioJ/STIatdgwXXSaSLJVUd25Ie9NSC+L8ZKEmbkkeDgYyUYLv9AE8cwX+KEB8JG
XQwxEbNcO3mZZpWD5f8CUkmg71yhttAGPtrP9p7P80aBNSaNKhsr0bR0OYr4vX2LQ/cYGRVLGU7B
qC1QfRZ6XClQ5HVw/bHfYPjXWaTQ3njQ03kEdgXMuSOvhF76jQGIXjRPl0lqe87tiBbaLTMoZbHs
omTgCTUJtu5p8yKjb6oysM0eiO3UWSPK15H5osqnYgNg5HFrRICbQcNDina/NItBMZJw1N/VqKBV
RNmntPGSLRHM+zNtr+zJza9wCk8mx5nuokHjibDkSQWQV4Hesspn7lbUSOB33GggF8+ZC8m90JvD
CiWQ289APQ+GwcMbCCven2s3DNx/br48YoGXUQV8lclMoD87q76fZXSZcWDGrAJ/RI++Ho6fJYJn
QBOZCMUF4hjqQSy1tg0TQUGvDIOpYws80L33GUKX0MsnpnVRmD03MOULiFDRGSHEde/T3Feex2aU
oYzf2fgEkPMI24XLyZY6Q1e9v8TpuMl7fWZUZe/IP4i3PzJmG6/EEUBAV6qrLD3dbd5Z9s+cifb5
gi1YPP27F8h30+yCEiYzcXrRGStuj/2TgCkG4FDcwNMaJTE39HCruCO9UhQIqc3Ee9iqDmArh5cA
VsxQ+beeehftTCFRS6XWl/Yk3cdHeFZdt8E9fEjy5q+1rKRJ99N/npFZBgok0vN9cnz5vCRgqSm2
yHuIY33WLV/z3JrvhQT0fuMrXc8PjgJYMouWfHcuflWr5hc7QXGngY6fPTz1Gv3rfdIQ2eht76S0
d3XrqL2f735D5N8WwVKp8MmftFsEmMyUXY4P8fm19vnMt2YOvcqJRBK1SglVpdRYwhAsQl1LbxrH
c1Fy9koZ59ejTZ6K9ZupZM5h7RlQnJ5+azaf/eDyhnenAhM6U64YGH4lLwMTZiWt/rAQK2qj2o+f
pqTJTIu9Wv648tw61fvoxRlN2X/Y1ond5tkfKstvI0N2055et9E7uvz3dp9BKPVrrY5Dn+3PIbBi
oANDNbXf/l2R/h27r9mDbnxdXrOZ/c5VMhEC6hfH2uH2wlShsKNqPTzWrvEE+mX94b0XMSHF0H8z
K4pcl9t80iC32KtvR8xZVHD/4UqNiFm0bnhNUovDn2Uizf+pMXOw2q6SFbICOufhoB/3lutMlq5u
MsjxH6+6S/I+gP0c0XpkuQH6VisqXSG5F9aBreIbmmzOkso5+HdHTFXniNEz0O1beQ4/1cVsoPXn
4+Dd9jwhB6+TgBdZwPOXF7oMpJ+um2zxp7dwxFBuJv6vCvqHUhbHIaIScgExXsU8gUgETUdEqJWb
VzUbknjFVK3SXM0l8OEZ3vgo2tBtoyg6KIwKbVCIsiteeE2N844erEkdbE0Jjwpq9i+qHQWuBoK/
EoR2fh6vUaVPbSXXs6JUEWfSUWkXwivfy/y+EDF4oqvZFsDUkRMphhBHRX5cnC+Smg+kdnX5XdxH
9sj07LJYYALlRZ2QnaIJNMYZUGmCQMCJNCITo0A0lE3Hx1E5Z+TJArvo3yQoPgqaoUfzXdvfhi/v
J9+xLWCKmDqyRH6392kBfmQfXWi0E+tszGIE5UoFVHo+ZRFLP3cOJvhDsSjdhClEZp2i9x4T5Toq
TSbIJnQhRfSsEGNYlhlNIF5eOdELHsva0h/o4zuGN5l8j99oU3s4A8yMq/ld5/q2u2xyWfiLPewQ
1x15Kpx/99tWc3k4YVQ57KfUJuV6SyYFVtkzVp6H9DS6rapLm2SeFJ/ORWJwz+vJD2kptYhh/Gni
a6zXqnndykHoZU/bKjjTnB0cnQ7W4EdShZEboADKwBGzh0xKSXaDp+KiiEf0Tc48Ey3M15fotdbf
9EsH6YCCNABAEH9ruhGO3qJ+Tmb/TMLYrhQXKBQBCiVvwZPo/pPFP1j0bYMkrzQy+VAMe0H1vBNy
8qgDGfpNw31gO9Uwn5j7lCuBSGE8m6Rv2bagl7qGjmsdMtPD7Gq2IKfOl2XdQhomax3WKA0fbowN
61GFUE5UjNyJ5/WtxjalSrqdPqkDG1O+GYzm/DYNLGvdW19kr2frPHFUqFiWZVjmWZAB+0EMZE5f
7TrglyVxLhyfSmcJb8w5rfZ+2neb1RXXowvhX9UrYcYZS2Yab+JGkN0U/qW7OzaoIGbSK7EQZgUo
J9hcRJHVOd49i5wUSdEhbx6AjZc0ZjH5zul6SMXEtDMfnxbU8/mIIHYSwWLcZXTBYN4JUl+WCqvU
nM/OqTKbhqmOq97iCB+dXmBdj2IGDpPZsjq8YfXTjlkPM8NkV+QSAJTfaWNW610ww3fUJR8F/cjm
8lUJ6xyytMt09XHra+uQmaaBjcngBumYEx0fFZ3Zf/7lLW1n/+M0nQoPJejOefTBF6HJkNTkkv+x
em/IIUIAKsFNR3I5I2i1a8W/n02q1s+Bmthq/6x1GeYb1OsF4QE3bd1C4gGx+nJuDc/lDdGAQpOd
x47eOQODHTSbLXiOEtDonYRdWjaVbRX5Qob/Cb+PstLZyP2hQev+6/flCgvzbCVROvUsCLrfHjfH
ZgI/1rsnMt4pxO53REnXmnMR2psF95528FCabB1XpTBQ+UAaAKsO8dEuYzGvSFS+fo6ItHkeE2DS
a+TtE4W8ccaI2WyCy04jxsvjD/Dsitnqj/4pMeAdZRm79GIfZieSJ93nfYVqA4UUfRR+CTgIZY3p
BMzN9h4506LrIGFJvgRCbtd8BPMX9mRTQrj4OXlgpICt1TLbsrW5RrBaT8/hgMZ6GEETFUyQA6nX
tJW/rO4S+EtcHGeNOHx3n1YZ4tJXonl0Tnr/HXOnfJroXUP0u8FdV3a+iyEcOWW7VRg4ypY6wSrG
ZH5iY8HDy6GMwI2pyiHrhLkyvLkYiT15kGQYvGnZRqPOQ9E6VsOuKAQK8eED3UExoh02lt18uHAv
f8Uf385n+yga9eGFTcBwicNGZlZasrtgFTwvdnl3+VpQ4m97AGmZC2p4z1q1IIKfJmwUPSPH8990
OOPnS4Chc3p0iRgCIXCbOGL7A43D3xSPP6WTbCSpy2KayosWpuR3iXuEYlXK20YEbW4zIuYxmRCJ
ggWe/CQU88Sq6X0w/5tRQEwPzpE2OuUySFJwqmi8QIvREoYmYU0XOlbdsoHSdActgolUzKeCmAGR
sgFCI+YPjeI6Kk38Engu1AHeF4yN4lrMjVMYssevHDMc5GCrvXNpQ1I7JMs82nS56ZgsE/lAG+TQ
XPepJ53bKjJ+Bu0EJ7FCiwsqhFV+bXbEmfk0qVBCXXQkZGNXLQqRTeDoOimQP1KX7X3LHssIFBm/
zZDbwuRqmPBpqdjU4JL1ndl0olVLdHIlgOsHw8AYNFJ840R3kQXGvdeFT1blfFur7a8X23FxxxIT
Z8gkeccVgMumJiTY7np20Wf72C3jf7JaBLNahg1zPmDe1iIcFLs3iUF3RywGi86KBtb3NjqtCJHE
qpDUE9GWnKdjj255TjnaD3IbUSiTIRiw92f+v+Nbhb4CqDTGflEEUpUbyGggT+1NCTs36+d/eCy4
25sdD3f15tcAo4X3epBvXF9tRBaY5P7Z0ViKylz0GyiRg0juP6FgQMZGWNRWCOATwLxffE1Svz+b
hqRREZOuetifleu/eS2VrmEfCGhhTE4cgmFKsgVsX2kfkRuqMKTmjb9O0UENPdpOuSabmXzRqnbC
j4oOUVNfdHFS9HXf3kONS8DvZnZEOWUeCwSScZ0EFhmNgWraXfCldx20Gq1pTLRwQHbyE3tmTyZK
Zry0f6+j5pEle0XwZpkTmPiM78+FzTopgBUUhZzU7jmQY4NT0MjxXhIfk4bt/AYgZwdU5F997Dlu
7MTbO1Q7SdTzKnstRgs/F7QRiaw9lZ0ZUPSRaFnDdVeaQmo+CVb2xSZkXYFkaakvnCsdj04sPghT
a7Xb7Fxd40XUhu/Q9ia/CwtvmGCTxF/kpM5FI6E8Hr+QNvb+quEr3f/x8T5HNrnMusH8+6lkiUDC
3Ukrb0rQjv02kH2f+WCmXS95Ba2/ilVHd/O4T+hTgy1SeCiArz/ZSM0V9P6jO5+Ef0DgG87a1YId
es00voDpPpj+hhto6iCGUn4ojsZK44U21m3vRRvfq97jEgRCD3Va1XG5GzltCFmxucz0u6nLJzNo
FP5NRT3QPepvrA5cVzPKeNadVOzByC/ft5/ULacOrzhYg2coq4CX7TEsk4T7olsBhEk74FCJGVQB
56xYM/RuPVb3bxl9WT2h417OsOz1we4qZscm+Z+vE4cOqJcQ3KhvGnj0BmrBnW5hpk02hRfnc60g
dsHhs9mmcV2Ran5cPTT6N9VT1TfFTyRlm+xvCAymIdxxGuWpziCuvLFExCTjBz8/xRmVbTr+3rNo
O/jHfl5Croo/2Hb3/LrMM/Uul3Rbiazfl9d58i/kGeh+uqwTc3zA29qcOit5ndVnJ40SjbOIxqgG
Ax36kLFH0e79e2WtpYIeB5iUrmo4pjq6KdYgGAt+8eH/FxD/A+6psNtNTnVu4BzaxJLRQesn+bEK
1Z8p9GxGL6z6E/MAVDPSJ4RYfSwkkfB0BjTTZO7JkiEbkC4uUGn0FB/MZZtWPouAFHgIAhPpj01g
/5tj2xVjtwRK9+Jh/akPdBvxWBwQ9VCYQ95fa8PXSLJlJIOLvK7h2zqP68qdoWde77hMvFCw7DNY
Skr9sazYdk8pFUg+dGQ3CFn/PVgqrJOGNKyjaG+8rTUlYcQ6XFxFcAu+Z25sYmPbYoZ1OCHmvEC7
AYReBvM4p20bmv1nGDY8mS+yQQLjFwWFeAQV/nLO0ddO
`protect end_protected
