��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR���[{�T���CK��TC,���:�
&��d!��]9�'D`�"9 S%�aQ�`!�6������V�W�l�a锦E(�\gC�slu�4U5=1�N�m��l�9ў��P���B�@+yg��=�}|֦���ָJ��M�g�=J�(:
5���,��Z7����\��e� ��y�״R�ߴ[,��V��ܬ?�CY/WAz�`̓�b8ow0D�a�0�>~���B<�c
�[T�u4'����ȏ��v��vw+����eErPB�vӖ��p7�Ew���g\k��&'=�d�N����O����Q�V���,?�㎴��1I~�Au��&��Fc���4w� �o|7[N���F~\H^���a�r�,��-ar�zp=���ҟ!�Q�|�C��W��˜HV*/�n�Py�7��[�1H�}�~W������V띱+y,%���r�f0S]j�/��~��V��P\��_ށH `�{����5����jB�=�N���cC�$��Q��D�S�c���ǹD���"���hʝ���m�m9� �TT̻#?���c��$�����h�Y�$�XBk��k����(50�_���nV��J(|+�H)e�4M=��]?U����64.�DW�8SV-���O��=_<��͹�'Ӈ�	
+� �|���A�+�9�:�����0�g /xw��S��:_.N���i(���h�q�t2�ٕ
�v�Q�eޱ՛I��e�]D^$m�c��b���M��t�V*�eܭ@΃���&]���<��F��`ڢ
��\�%1`�ꆊ�*L$.�JYpw u����Ŧ_�jO��J=��X��:�� {!+l���+�-�N#���7��G]��Nk�Cl7P�S⓭-����z?��[�aL������EKg�U�RƯP�����̇��ڞ��o�M��<`���W��T	�_��b-�-��9e��?�`%J�d��^ay���x��4�$:<?|��,�&?���I��i�%��vU���ZǣP�jh�#�ؑ,�j,��RK��j���^W�8d�B.'g� �#�Y&�A6�
�5�J|�"V��1��a[c�0+���6�*{�f���/ʊ�#XP�����%����VJ�.������c)�}"�M|�'�����ی�����w.��j��� ux=�;���������ڐ =pCx@	]"u��o�{��U<F� yA�]����E��L��b��P�@�2@�>I�st�1:R8z�a�t��,Ek3����N�N�R(�����`���U
��7���Z���t6
:Z���m7D�L]�A����}ٌ�ʙbu�S\!V�_���l�$��*>"�B�L���`S���A#Dn�O�S)�c�^Fg�t}��^�r�T�C�c
1pC�#�V��NYV.�*�7�ÂB6�G�wA�Ȓ�Dงտ�����S3���K�0�����Z	�v��V �"Tt�m+�U��%a9)�[G	������1<���[���v�m�	�fKHޡR�z(�6�i�H+\����$/�*ն	�2Y@�d�/!��~/
 ��z�N������;�M-B0P	�4��E[c)U�\�4�2@�b��\J=~��̞����)ߢ���2�Ρd�jv�)���0��:�
�� {:�� �c�x���Q���~':�x�n����']u�B14����1z�l�<��rgwx��t w�ғ���7T%N�Bɤ��ԫ����@�3H����ᶪWZ��^�O���ٻQw�흣}�fkf\
�8Lh"W�rC>N�r�������eQ���F��+�k �L���T��H���W9��8$���ƽ�4�j,�&��.S����4�^��'���O�ct��.|��Z��l~���P�X7z~�|�Q0��p"�.�U��l��*X�{����K�wx��H��l�ؗ��$���O���p��	X򲍎x^��ܜ䙯��N=JKI<נX
jȭ�n5ʦG��4���<簸�(��D���!��*�(^{3�����~���)8m�r|/#鷑/�s2���2������Օ!�Zɾ�7�����!I�r���FxZ�@�o� *��e�~/��,��svLT{��9�)AG��gg�hJ�柯8­t۶z���`oYM�̅d`/��<�ٸ{�JN3<�k"�{}3s$X�!�è^Ԣ|�K���dV��2�Xtx��>�b  {��;�M���U��/z(�Y�_�K��x�p�BB��t���|�r�=�<�pM���~�T�������1VQ��lLg���R���+�L{� #�>!�t���Qk����D��C�{��M�{�D���E�%I��=L�H�0@<�lC�9S����,�}��~�;����O
�ɪDԿV�`���/����w���#N��&�1��h��	p��T٭�Q�,�M��:�]̫���xQY�%�MwijjQ��,�#fT(�L?[K��f�$�l��.ہ�j>�����q�o�̥�?��L��l��r��j�W�+�Pa��#%E��p�,��&���s��s|��E���U��%}=[�pñ�#�D�fX��M��%o�w&�5[$�7��	��;��.p�GoRОʼ��X	�����)B$�.ₐ밬Y�����HA���VC�����B]PV��Md{t��tH6�9��0-����!H+�.��y��:a;
"��y����R&�ћl�|��2�"�hi���6����"D�+������#��>ố/A����Ɓ~G$p㗜~2���#@�a�_��q@��d�Y��̯�@hD�Ua���yuAP#}~�,���j���/pӣ-d"���{�xV�h��Z) ��͸�fI���R��In��i�S!��NX��Jq1rm^�bY��+L�}ṱNz����]K�����c�E���6A���Z�{�c�tl/3�B�� ��i���Z3�¶@ls�A�AB�R��$��?�cdΞ%��OP� ��$D�֟Ť��9��"^������mٶ/� �g�<�Q|Ӹs�l� Q�\ %�G�gp�?�������30^�0}��;ֽ ����P�����_W������^�]���˲���z��n��%�aY�,��U�|�"���7�Om�[�_,��(8ߗ�!;Q�.�=�I��h���KM48�Zibޕ�˾0�|�GrG莋e��lJ��堢a�u5�0J�ǽ}'Nà���N5�"��l��3L�/�!����(q�fZ��j ��ɇ����n�Ki�nY���7�!ܟ����-3N3-���4?\vx�,x�����>~�;k�*c�-���U1��W�A�;|{����OV,R���=�vۙ�!B�n��V�'�1���"-�a��"�M�YA+?�u���:� ��9I�}Y�j�XO��I�7�����Q�y�p�k}h� �V��m�=G����U��u�ϣC��|��q�r��}�m�5��SĞ��L�u�� Q��"���B!6Y_�9<�Hg��� Dr���盓tC3,̟Ms�1�������1��Ə��"�u��\4&�
�z�+L�_�:�k&|�;6ٴ6��Beg�4��A�-�EY�����6PL �Cp�	5�e���v���mC�x)Lp���9�y�p�)7[�;Z�����\��dT�ΆQ.ǣ/�:}�vc��@z=�v#�-Hyq�(<�"��P��L�V�ƫ����	2+Ho�\�cI�b��4&l$\#]���F{E�����pbø�;�I�	�8Ŝ4Ԧ0�S7z�K����fU������	(Y��$\Z�4}���xV.��5�J>`��m����!���0�̣�"�|�v��|>���i��XΛ� �@HA֊��w ��n̂��~* �X�Ϯ8mea����q��g����8�ʈ!� kT���W���â��I���V�_h��j�K���,
� ��H���ͯW"Md����qk]�����,\C!߸�a��hU �t �a%�,E�.�F0�־䡟�Tw���
K�@\B���;<$��V����R�0��	����E�2R����/[��:�2�!��spE�rk+!:���,�խ~��1�a��LF�H�+br�י��a>>#�BX힫]���S�����d��pq/u�[�����m�-.�o������02W���Y����}?�#��
G� ���^&���e���3�m�S�a���І�Zh�(߿j��d�����,��L1�\��=���f1���sP�׽[�z>Ĉ�����jȥ����|]-��?_u��ˏЎK T�0I#K�Hܶ��Ћ�q����?�n��2̫�"���ο�*��>����F����u�]h�z0#uV�`a���`w4����K@ޮ~������(0U��iX������^��+g���Ek/�%iq�[~�:�%�U�F��Aeτ<�Ѯ���b����@K������9¿�ޜ��\/�ihIϿ�_����=� �k(}�?2�����N2 �4�ː����g��Yp�|c�2����j���jy�' ���1\��^�{�$p5��nbK��C�ãrn�⸢��dK��G��o�Q��d�'H	*%����w�,�3�3"M�ps�Ne��pj[$jl!;�{o�~�P?�]�tq��\�]PZQ���D{ϊ�\���@�dT+���]o3H���<��I�@x-| ���9<�v��8�Dw�$_�S"Bx�����=dG��R�h��{ᆥ��#�~��x���`܍n�R�~yu��p�Zj�.���Z��H��,f����3�Rl�3�M,1a�b}�9�G��Nt�%�"������P�k���r�"LY�9	#����d�q�	�;�v����>��9��;0A�L^M�u5:�\��ԗx�	Q+ �*�w ��Ji�%�c����!�/����[:�l� �E��izX+ݴݩ5x�h�����l�U.�Û�;	H�3���ۡ!��&
�_,��1����:���y��)kL��+Z����Ɩ�8t�H��	�n����	%Ez�C��H��I�x5<#�86S% ]:�s7�����ba�O��"�8�^Z�O��T��v�ޝO�t��{w��f�_y1݊�'���ζ|)���-�����?-�/{�y�
�'��P[��E�%�>A�]_���%�����Z�m{�Yk�\t�T��˂�����fW��j��G�(J�q�о[ Тh|j|۴k�V�u6;��m�F7��\��?x��/_FP�U�_�^ۓ�G�]�rA>�H��,Z�8��}{mE�D�܆�Y�a����u|�=���(hd?��YjƇ�sE�s2eu^��Jꯅ�o�(GD)�4�^8TK8�2b��	�W��뛥�kd���y�,�4��!�js�^fQd��[��쯤���!�n��� ��a��D�L�	%��wL�Z����F��/����˷c�� 1b��?C	̧��W����)g��^��,gު�f�0Yt,�Q���qW9�x��I,:���k��b���r�zfPa/64��'��NEj8�MR���j�� ��I�+�L[_sw5�j�v6�L�a�*�]bz��4��z���GOg�U�c���3�����5���rr�`��ph�'(��~��2d�Ղpl��%��2Fo�"g����I����A̠�ey�(`��t��Q�)j�(���D�=N�^���*T[b{��4+�Ä9�ZVe"M+����u	���g��0?�n���f��,x�B�Il�!����J�lG���)@��&Ve�CY;�������%��^�j·�����?�����������\m������h¢�+L�~gâQ�J��RA�q>��Z6a���*�#��x�W��G�_���7y���y&���CZx�b���0��a�CcE��f�Ye�ִx�)L�@��_��c��ו�m��F�!�7屖`��9�"�)�hE�ږ)�j�_��9ɞ�
8��(l8�tVr@dd�=��	����._.�1����P�<�I��+���6��$��"��!	��Z���r��v�Yq�!��X\6WVR�W[eQ��Ԏև�s���͎�8ۃ�v3�3e��-�.vN�upi�I#_�Թ��W�+W@b��NG�2P�V��KC�>�t��)��k�'a�KN��b�Z4��)�����r��<io���Vp4Qaw������D��_��*:��ѵ\�/۩�D*O^�]Y�^�*��u-G�}� 箎e����l�Ь���3��`����"����դ[���{����
>X.#]7�{k^�����-Í�� �:�=D��B����ĝ܋��aZm�]���+[�/�Ɵ�[�`����Nw��}����(�GaQ6���"^~L�#w��jXYub�0%OAu�B���(�LI��ili=el�����S'��}�i�4=^˵,"t(�`h����+b��$Zָ����)�k߾�5���H|F�9��4����K��Zs�ɨB+�KZ ��؀���	\NL(��cW�Ws�?�b�T�t�/�-j����r�� �<�\�9��qBص�^1�����Iq�3#�AQk�M�(�G���kՐ�1���$(֎`S1���]��/m���)a2�K�liXx��]�@���#���S��S;���i��W��u^DD&���z�C���ֈ�a��1�3aɧ3U�F%G����)���K��rw�[���¯��s�V�/�# �\<\˪�l��q����J>"�"ľ�#��2�+�� �����#K�H�
��F�)U��:!;���V~bmUӇʆ]慞Ѷ:��V��lr�+��"�Nl�T�AQf�o/��%�Cu��vOn&�W��}���1 !�79 �A� �8���E���%�D���˥�_�K4M�:��6�`nm;��;�CW��M�h�l���Ǖ�Q�Yۣ>��4s@I�t�0�ߣ��I-P������~8�T����^(�Cil]���=	�zB�?�2f������y�K,0oW�klT)�r�����Y+L��$Z6�q�iX��.�9߆�hޒ�~�kC݆��&��N�HͱC�~80�A^�r��V����,E�q��'!����@F����vVr���E�{C��;�Iɐ=�ep��#á����A��h7;Nd:C���S\xץu�)�˭�:�fj��I�^W�t���Obצ���BN� �8�b{ә����n4�=�g.�	4^�b�QvA��)�K(�ޫ�~~�(G��'A�R������e|��[��ae�̄Rў��k
����<y~��c�p:	�{�<�j��L�*/4c_��pp�A��h)H����nK(�zY�C��v���j��QD7Ckե��ʮ,�E��X� �	R&t�$Hr��~w�vOڙ��NWݾɜ�4q��ŇA)N&����.�O���l�$��nI~`RR=E�J:k��Z�
QO=���	m���Bv�Y��V�k���y@��.'����H�	�wWws�!���W�Nk�Dt���� ?��bf�>���o3T���܏_US� iX ��]&��$��kC��f}���O����s�)h�<C �Q��*�$J��L5����F��B`�?X�a�>������6X>[��u�r�v��R���H�)���Ӏ�^u?x4+چ�B���:s�� ���.��ǒ<J+Ϯ�,q���j��U?Ф��ttxWR<>
���qi=`�}��rmؤ���Sɋ���:����iT��&8��4��n��=
��"�0�?� dx" 蝗dˊ���O��9�T�=�gl4fS�c���X���av�������e&�`�T���\��s�qō/{?���Ac�ϰqo� �a�ӏ�_g=�z����_�g1���v�|kIo#��u�F��ԬC�b��_���'�M��C�~l����
��iT�t�Ҕ����$0�x�Q4B�,)��Q����^�vd
��(��-Q:b�	A�v�C]�cQ�����r�{���~�_����I��BQ�yO�m�/kc�c��,�X��?���i�5�D5��T_pY��R:���ʛ\V\���7��o��o�!%�&:dJC~��X�<�J��n�`,�Iw��d�����O��"۰�����H�[�3C"�Ϥ�K
�\�n����H��*����w�������0�%:"2�Ǝ?*&���4��[a�`�s�}(��f	g
	��`g� Y�@3�����w�SI���%YX�@	����ɩF��q��7<l�.q�O��<8���u�x���N���=�*���9@ax4��{0_ �I�/G��)���:�i]L���c���`ns4�xl>�vn0��N��S^��lSk�r>��^bn�	T��	.��F��\	}�"���S���1���M�R����B��;'�>��L�����}׭�_4�Z,1�{��π`��ґ�J"5OE����c%y����a��N�=ś�r=a�r�1b\"{+�9�-����D�l��@o/�0���[\��>�����
ַE�[����E����������kh��)N�T9�N�мf7�}8�����V�;�U�����PM�7Eo���:[ՠxPS{1/n*\�ޥ��?�#��zS$"��dE����qr�즩yEάy������dS����z�0�Q�9W	�\�f��ԙ�}�tv@N>z�3��L�6�va�6�g�Ie��T��l����|Y�U@�S���h](N6�t��9�v�:�Զ���O�(�+j���)l��\��c;.��]�F����}^��6���(P|�#~�;���m7 /K�ڍ�ˆ�C�6'�{�[nṕ]� E�N���D�C�&C���"U*�����B>�2x��6��b��F��L?qʶ��&�3�ߖ��%���Wxk�}֮���f���R���E���/��l�y�.�,T�[wˍ�Sa ��]̿<G���v֖N� ���ۻ؆?�b�f�DW��b_�7���LKC��F�W����xK�o�u-��(.erm�S�蓟������tm�r���wl�aE+�s����H�>��P]��p��e��/�&��Mf^�I�-�C���_���-��}y�
�[h�&����1�!^r�)NB/���":]Ҹ
��8B�� ��k('*�%�E۠�v��j^�G���3�N2�u�\%�4\���4zL�$zu����b�! ��A�4��T�x�=��R�E �n2n�l�,�9�f��:��[�D�d�0����g���I�$u�KĬL��D(�s社9B�l��~B��b�PO�p�,gjk/�{/�L>_-f�Dp�)�x��*�C�U����F*��~F�8��t��\hאvT]�&��Ě����Q��%�$��E(��T�%ʓQ嗄��<���u��;��6�[g�M��
�HQz��@J�����؏���<*y�?�m��1��!5fJ4ស����of��'��g9��}���*\Z�I�b6�T"��b�=s�
٤Qng"�1J2�
-D!Ga���Y'���F��I�$
�>σ��ב[�睑WQz���Fd��٤Q&��}n���7j���+P!��T��I�0�Z'RAl����Ծ��#��kq���k֦2*F��$r����v�P�!��K���}0Ł�F�&��O��B����_;�I��ٓ��*�4��t0|h�y�A�}|[��
�`�,9b}��$��~q��$����	���F�lk�:p��䟨t�vp� pFz�f���pkp�ˡ�w'�l�s(.��'��ߩk)ԔI!��%D�;�	f�y�� � PlCm���_Z�l;���oN����`��Ѓ�m�mQ[��;د�?���YT�HH������݉�6���Ɇ���
w�A3�^���M���E���. A.�$�l�g�)���'tB�\��(o��K�$.B���@2x4�L���Ll���vl�Uu�}O=s�z��?|)t�1D&��V�� �Yn���B�_\Y"4��n.��� _��[C��47U�J��*hcH�v�)L

eX����k'eP�w�F*)}k
f�bj��o��B�G���ρ[bVW�0���dl؂��O�]��V��>Z�ƘY
��w�b�p쪅�7����"Sr�<*|/[Qs1B&e7��3��0a��(��r�!O�Y$6�#o��!Ias�cd�^Ŋ?�S��Ҕ�$W6f".����#��  6x���76) p�jD�����]��q s��@ðn�L��YN��U��e	Z���3PWo�tℛ�4�� ����Z�c�_/"�=*�j�)����l�w�*0�z��l+�Ȭ�YqY���Wim�u		ߦ������ƄK�؇ {�f�(�F�zp����>�
?��u����vj�
��"�²�Ɵ����P8��\�e�7<u맔�	��'����+]!��A�ğ�`��cnYf�zg�qH5�9J$�b��T�
�d�Ff_=����<�&'�YQ��ƶ�	w��ݓ�׀$����P���/�>�֥Iqj(���7܈��Q)4�Y��7�ex=��� � ���qo@��#[�CQ6�B��K���%���9��v�c�`6j��,u1�=O����s=2H���i�m��Mؚr�a}�B�;+�3��,�a�D��z<��O�{-�L�(cY8Իlf��M�h�E٧��~�.H�@*+TrH5�����*@��T�/^50Џm�Ŗs�d_~�|��h�Jqu�}�S*۬ 3z�ۊyQ#p�%?�M�ůWf�ue���',솚-�X�R:63�&�����ͥ=̚os�X)Q��V�8��oݥ�	�}�\�3'Yʸ\�Wg���>�������>&��di/2��>�F�e��D�d��,� ��1���pt�@�H�]i/�	T�N�\�zٜH9�X5ҹ/���p_���z�ʄ�'�҂�p��G葯Ӻ.F��sB���ƅF��-6�p��NQ�Lz�zueѯ>�!lĽuW�=�+}j���.�����D����YJhFb�"<a.�W������^�^�33�-W�3qA�'Z��V�ߒL.����L�r&���K�f���.9�m.^�Z�q�گ��&��$#,u��
ku���A{���C�W���j��v_��AL�F���gA�fGӓa���c�T�`fE�s6'6�~�Ȉa;\8��Z@cW�� ��)��/�:���ڼ3�sƪnB2�[d��N7>Ӣ�/o����
g��`�,����n�A3�㷏CX!�B&�!^PP��#-k*5P.�|� "�K|㋪��h=,]�.�t	d�@ɢ�Q)�Q�9aw5�>�F��.;AH�Z�wOm�l��P�K��AjI�x�#�y��[�F*��>Ɨ�dl����)x����۫��{A ��~|�'�1�^��=px/Y�Hr�CKU��~'�ޕ����W���HE1g�&W���#�T����ic+j!*�Fyϵ���oX5�!Q�Ţ�o �"������1M����)ͳ��&��oc����es���MQ���Y�tX�zZZ����AY<�s�ȁ�d[�I�v������^�e������8��"�X�.����k��+D��z��r���)���:n���L�|��y6O�UTw �mR�@7Bk�.��J�:�-2��Mq����?��jN��sO�t��}��g�5%Ҡ5B@(��Y��X&~"���1XE۞�9y����$x�nz?��
B��E��oeݗ��n��2K���d���#����B��G��#�/�t�qu���.e�[�FE3o���ˍ�Ú��9b��%�bʃ=��j�R���7D!��i� �)G�b�Ӵ�<-�w�X��,����ӛ�O3�n�JõC{��O?�O��6���A��59�2 ;i���;(���ze*~)�}%���1�������eNO�"�%���U�<���n�o��6^2�ƲY�{������1s��B�>-��e㨓f����馿�&���O!���S��qc�B���)g��Bg���ct�tby�����,8�KEP���f� ���ZU���p��RZ�<�[#e~BYj�Z�*���tI��&N�!��lP��=)�c�ﯼ�/^#�5Ϣ�!�Wōǡ�i�������a:�?$d4���7��7HU�z�ey�,%��^r���ί4����x��p�bO3���.l�b�W�mȡ��	/���L�Ȑ�Qj�d|��x��̀��C>{Z/��U���Ǘcsc���X�;�r�n�4%��Y�M�7����8-1�,*SF>�W������Ea]�k�9�G����t����o%)�]��=d���M�e���`/���x�c���bS>�N�9�r����x<<���`����o"D�ͦ�g"�:�(��)s]ÁE�9sS@�(	b���"�A$[�_5Q������yW���s���c�������J�?�����"n���\C�ܯn� �L;���$���~�I. �bD/R�Fx0�U�,J#_)D����\��uJמ��|1&w�'b�R�m�[���V@6 N�����(`m!�qQ��d��R鿡��
�	�q�*�\�>�g,�т��iw����2����0柩Hs��4 i"@�Hi�k���j��,y����Ds_��T��y�E
�͵�:R�vU*[�X��FQݎ��POo�n���uF��s�[��``�����=J�M_�*��IDAe�M��/B���FqV2FnX���Zp&@ =O�c���H[Ud�P�}s�G<�90b��}��s#:����*��1
��
4_# a�W,B�<(����L�	�?Q��˼$��#��h��d>�U:���o}��x��B*d>���D���F��@���ZZ�c�;p�:�p8�ڑk�	8g,` \iF�E�4�J;�![N���8��5�e����1wen;�_XF�b7�Y��<��V��Nm�BZZ����c6�`|u�q�ʶ9�Z��N��v�.�
@Ι�h=�H[XG���'�Ҫ���
��b���B��Y�7[mf�|�G�㷢��s����q��oR$��=}GE�S�]�RTm��x &%�ra+\�B�h�,�>C�8�s��
/�}xO3���ZH�u��d��ԣ�}�2���B'mc�7 a�نg�mF��ѰySNI.h.����̰���Dd%��a�j]/V���FmR��d8l���u�1pYř���@�w�Գ������66�\::{t��Cp}S�޿��=y��p�c���p!7�U�S�Ű8I���k������D4����'�	�NE�a��t���*ť�4��XO�$;�Y�ql	��ܻ���lx�ú�)o\5�+A�T�T.`�sO^�W���j�ЫM�7�(�溎�e�N^vͯ<W�舚IH�n��u�$fփ���oY���SDɑ��`f�y&�8��qL˄��C:�$J8�(����ʤ�e�3y�7x	�Ӑ��߉C��9Ƚ�p�U�B�mP�0���s�pa�=>DW�\�a-ͮ�6�u��u^��*Ƽ�w���Z#�9��/ҌJ8�:B3��j��ƍ���{��:z|8��F1�'�$
�ф���]2˷���Ho�& �$*Ɣ��sT��=Mr6u��^�c	�E��GB�*�z%�F�Qײ���K5h�n7��qe�p/_U�_~M��r�<��=��g�%1��ŉ���t���ѕŸ(�dZg���c�����I2j'�e�*a�5��;���A3�?Tح!��G��)R�@0|�<�<�	�U+:O�57�6�8����چn�*U��-�,����]�*D�k�I�|t%Su"6u��Fr�h���G8*H5����4�|�es>��<g�2b�1}\`��r�Q,t� �%fL�+���>�U�ip�_W]G:��LK����(�{�픚W"���dra��l��x�U�J�Ic\�o#ۊ�E[_��@	W��-m�����S
dE`n��]X�6K�/f�	�H}b	ȱjb�߄7��'m
0�*#�e�_��хm�(R����zM�55+
�̱��qł��W���'i*g~?��#S�j�K�P�k5j����������@︄��۠�F�r��ka�f�(eh�^Ԑ�l���F���ӥ�t��)�V��X ����}Z�U�z��<X�\M���J�k�m;�VS�q���?�EH^�w��~e~���L�q��j�,'hH���8_��� ��8[�Ó�SϾr��87�\_�y��Hy���1D�����$���M~_�Gh���P�|���7�~}jO�"Eԍ���F����kxZ$�2f�sIzgV%!ͽ�q������l�fJ��%�u8�R�����6	BEå�iг9����%*z��Eٔ$�\���2PZp��5���@��9��~s��$�����m��%��*ɧ
�w�`XDs�@I��YU���x��3�K{(�.�K^h��d�ܖډgʕ��3�fH3lG��~�䅝،�@\��Mv�1|��l�"�|wT^�����d���
E�-�"T�j4�C�'2^�O����S�_��Wj?��(Ձ`�G���L~w����ݞ��d�>�?���.d-04 4��y��+��E4e�g>9+$5�`m ��%���w)�7(\T|Wd=5�JP�������e�����ۧ�+�߹
���Y|q^����&��_β���
h#sxX%lJ>�9z�����R�d�'�E}ji�(\nCO��H���By��;����~���v!�<�|� �T�����/���K�PG���)��_�(C,�̵p)H)�d"{_�sS�Ė{�"R�^=t�;�N@3�'��3�A��w�,���t��o�X�Y	��Bį�0ح�rq��)n�^���ż����V c8��Yb�|n�'�i���&��S����N&��(���|���O��+�rx�u�9]b���|���ΌF���Y�j����M밙��׏!���5�����J��s�f������-h"v��9��Ռɕ�ã]����p}��"�KA�P'���0�O�GP�c�{o��c�8
����9t�*�/};���O- �� 2���A=I���~ZU�<^��>$zM�䚞l	�;�:�ĔV~f��3Dۆ ���s�톋V��Ŋ��r��OrZ|jQ��� ���d?�08�E�t��]#K����P�(F��!oby�WpI��r�c8�My��,[9��$	W2K�\�@���XR{(��/9�n�g8#�.�2���Z��ie�NBT�."��d���G̼0���)����F@;�.�Q��.❼�v��	�6��
wjrR����d��)-0o�mL`j�L|�>�lX8��
�g򽡹��@�*OKerGp�|0N��P��d��F�5�RǁXJ-��[2��|���ZXL�,R��\lXink��C��s���ݓ�?<�N����J$ O� ���rY��|���B�s.���gO�Nb.~g!��Vu����G� �f�c�{F���P��o�L9'�d@K��~�$��i�y�����-B��I`ݞ�2(�r�����%�jլZ�=����)��t��a���,������eo�"K@�,1Z]����V�*�?��!�8i�&GNJ/��, ���mSHF�ݝ���O�-ܗ��r���EDYȞ�Df7)_�GD�j�oS+\mDE$���2��.�1��/]�2Ǆ�5����&2͇{;�-k�e|N�I���NE+B�#Q���<���6����6�д������RN {w8�*��:e>�AJnh:+:� ]���4l���0(jz�!���6Q)��p�qYT�6�z�-�	�GA��j�������P�Wc>&�f� ������c0/��H|�頲��z.f>!?���|��tp>��y�'2\c�4;�o�"�r:��mB�9s�|��ys
�My�����$�ݽp᫑�K�������u���Y��%n]k:䖫�X�_R��sƈ,�g�8��1'���u�t�F��^W���QB)�*����,��ϑeP�LItH0�ƌ<L��(��C�涺��!�|�ޯ9D������1[��P��Ԥ6b.�P��v�H��2b�͌�b��.!Z�P����l�Z9D��ϩ#g�;Ǐ��7I�π��M]�5K�
���A�;� �4���>}�$��u�?�t�o�H�?���xӍ_c&��򏿉r	��?���4��Tĉ#<Ep"�y��ؤ�ƭ��4��^�����2UW�R|���]�ȝ��޼ �B��o�y3]x~||v��4���>NÓeJԞ�v"#T�o�Ye�1[0�Ʊ��N���L�m�\���0Ztw��k��㟶�>�(]�^Ӝ�;���j�Nv� �B1u�>�@�K�$��"��w��M��$Ρ8V�ɶwй1J�J���{5#���rG\�AI�T8��P���K������w��e��������{�*�G⫻c��o�8�CF���&f�a�Y�[��qx�3l@rU{��L�u��4�2�JL7��v��j&+q� s߰��#\��>`�kX����4dNH�
j�|�r��pOKn������f��� j���Y�.�ְw�:��,���JQ�A7��<����%�砯,w�9�����(��=i�g:�u"���+�1UBI��4�<K���i��z�w�Q�ܮ���Y�a�ЬΜ�:&e���]6\���uN��H��2�� 0� �~-��]�'@"��ra��%u���0<ڷߌ����eOQ?��(:(���G���~��	�ap��_���޷�ߣ�t^p, ���A�]�,�d_%z���g�|4�Mp�g��&+���V�md�����yP�B�D��;|p��C&��M��h���N�1w�D�.2Mv�k���!�}�i)�Q��s��{�S����.Ir��.Bg��!�L�����J�@�m@�&�M0THb��Њ˷��7��/.A��#�(qDX��Q������c0t���V���Dx�.GfA�'��B:�l"1��3�z����O�H�4��Z��7��;��_KڭDVU� 6�����e��p�ĩ���n�5<˘&_�jv[�=�����xM��zifS���T�#o[��'���C��F���CM���J;���?�G�)ƹ4������ȱ.��c�T�vz�^9D9����d`g�XMg�IRo��@m(Oά��)�%p�Q�ׇ"���ҷ5�*�Tf
�֤�b�aw�whi�^xޚ�C,ߖG}�7�2{��$ ki�Q��Y��Jդ쎺�J�&y1D_�C��~
L�^�6%���=@ΙS�q\<S@`�BN���=�t�n��&�a2�����Uw�+#�nH�3c�!\
�m���R��?���GY:���B^��zA�!���ܫ%�6���L춚���o�d�e>���V}���c��s�f���c�AΒ�VÁX(��Y�}��@l�s�q#��*�����xk�VY���G���w�}�w�l�rRyIC�\DC6���  z��k!_Q��j5�H�y咥�D+�{�Co���9F������������G3�Z�SH}�Rv��BjM��耦�s.>�#*�-�����뤙����Ra�]��!{?F��/�6t{��� ��9��GS}vE�s&�=�}���g���*�3���OV�w�mۻ�[��`f%g����"1hdWZ�Sp�������F��^~�:�ܵ���Ƞ;����#�B�v��F���WY����|!>�|�ǡ���nu�v ��8�0/0�MT����?GJa��+�F�����$)��ф�#�-�PnL�B%��;�i\S���C#%
�㰆�}�z"����W���_G��C��F\'�4���B�)�	+���<n�8OF�-�Mkr�҄��v߷@O	-�	v�@���z)Hy�ϹT�	�_N e03R��C14��p�R7Io~旓�as���2w��<'�#�a����)؆93:2�¼ƿ+g:2� ��;J�ݽú��9-j���@��27���)���+��+)m�KC#M�9b�c�J~�+'-�hg��Da���-Tƪs���f����x$�]�� bUX��n$q�X��*��3Z�5�R�?_�
���ٛ��Sw̢Ő�.7	�J�D�p�sw4i��f�>@���QS�-��7��+q3�)�W��}V��Vdf�G�1�8�̄U^�2�w��'���ʡ�gkB�'ϴ�q�>�l�,��+k����~(kC�����'��-�@ͺ��l3��yV	�9��*�&��R?/p2N`{�<Q2�F�Yl*���2d���4i���K0��W�r_�"j|f�z0�1�+I���q�~�j9�zm@B�z�3D#X�������7U�;^$@�øv�?���/�-�s�0_�w2�V��E��?'חOԴ̎��|��Ǡ��1�<�I�K�	��vl�Pj���3����©0�˩��0:�V�<ݏJ��p��-�ږ�..���nG!�L���qy�/դ������%���5���e:
���":9�(Y�s0!�_�4|2�(���HJP?���p�E���K ��Ȩ���~�8*�NC��Qp���`X()�±���Ǯ��z���I���!�b3����$���+�z�#m����.|Zm��뉻���i�Z�f�kc�ꬂ�,5�XZ��H����V{���_��/	�m�Rd�_��Ғ|���/ʋrpil����'�Ï��!5A���H�cEN 4`�kU��J$(s�e�<v���������X����[��-��Fr%�O�X�&?��e�{8:��8GU:H��De�;j��A�4k���	6 _޷PHm��Gd��= �0��/k0P��$�����ׅ��_v.�ǟH�+a�;�օl��S/��W�x?�0��O�mw�*e���TL�9l̫q�����8�,g��~�ֳ��I�����P_�6�t'�uAm��,�8��RyX�"Rܯ�.:���7DKr�/��0�_S_��-2b����ҔFO&B��5�Y��v���H��x�YٷWd� ���8�cq�Z�ԇkl��t�eI�Ly\��"��^u�%lw��s����15���4go��1���'}Q�,j`�I��2�X4I��D!q0%���F[����6L���:(wT�Ǘ�y-E���V5ei�F���0�Wj�3?�����9��>��V�1�����
@�\�2���N��yMr�ƿ���%�?�����< ��w�y8���u������Ax�M�Ύ�/���vPŎ:�V==�L�\��3i��� �ZeRX�}�uxڋS�.P E��
�Wަ}+@6|�!��`�|c={��,^��B������@���g�3!�7��������P�6��G�Ӭieqg�f�&$
��<O��N�h�Ӣ���oX�Э�Q��C������l[��}�'T���d����j<��w���� ����*�_�:�bK�ろ�ҡ
'zC6�f�h'�pP�t���?G�5�n���[I�0���O�nM�5�< +�ѩ4֕�
p5�kHdJҠ����6�U.���q|F/����S�L�=��K*(�Ġ�5�^�Wl~��t���Jk[]���~Jl��sԓKI��d�"��w��\�6���d$\\l���美.W?(=�p��j#]�������#gӛ�^
{��;��}�Iv�v_V�˾�\�@s� �����S�>)i�欅N�X��~��u�=Ǎ���b�Q���
r,s��7BI��e�;����d��X>�Q���*�,{T�&���5�0��
z�M�֥Q�HT�AC׉]ԭ���Jp���1�4~�M�'���D���<���z�7H`V��o&�����{u�pP����c>�F@�_ͺ�KouȮ�($��W������]C��I����� ��JN*�`\,F����G�ζ��6��c�Yv�n:�����	����,�Ńm8��v}r��K[O���4/��3�R`�$|2��W]���A��=�:��3#RL��;g����]�r��?���~ �O�F��r�ä���~eEə�n53�#p �FW<l� �?�u	F�*��`Q�����f�J̐����񧩡i�Bˍ&�D�@��%����fw�K�6+^%��c]�Z��87�}���nhrH&�c��{S������S �	���ן�"�I��O������'2~��_/vc���K+�~�Y�N!��[	^7� ����:9b�RK%Q����~���y���b.���!� XR�=΁��)_��x:\&���Ldl8f��!g�ף-8�_����8N�8[���3��<'H�� �<3mV2Od,;�X]`�����.׸��!�8Y�Ԫ�g�� ѷ�ʊ�\գ�ׄ�U��I6[߽��}��(������Ӈ�;h�
a�����3X$��YZ��7n�lc������i�畘VS	���ǲ�g��f�����\H �o�_��=T{:�l[=e�T0�S������.9�����7�S�L~U�1�Z���p3A��{kK��t��3+I�En�j�P���g\H}�M�i�����sF[��Ɖk�
�p��+�q�'enO��-P�(}���ՁIR�� %4��*�a����r]w����w�$J�UiZo�"h�,�[�J���qGo����Py�ܿɹ���O:N`��?��*�t����e�j��$� ]D�e���rd���T�HuL"�m�x��ڃ6��_Pi�GSsYng�>g|��1\�	)��"�b%"��&�P�P�՛?����ZM�1K)��E�粿�|�9?�p�I�)��>��V��5�
���s�dMQz|���0P*��`��:&(4$A�U`(��Ƭ)�ˀ�2:Ÿ�\�ͨQ!��p�����]�E����ڢ�B5����3��$��?�f�C��u)sa�����FB8q�X�� ��!�"���p �@7� �B#��!�� iON}(?����.�x��{e̝^�0�LIf� -��� �avOC��?۾�A�'�H�{�q*�g����џ��뷡����z)�.�5��O;�9�y1�p�|��o�__��t���^'��}�|�qBL�J9��f����m�.n#{�5�en��`�n)��_g�ڱ��iQy�A�O[�z���n\=b�%��J��@�@�[֓ãۜ�q'��D�:�I]n��1O�b7����z�����6<�?B��Za�wXڨ����c�K����g�{��M;Ԣ�V�;/�l�ǽ$	7��٤���wL�a�$�j|���ݶ��#�������M��y\i�A��7��5L���b�p005(�X�K'!�@��ڭ�3�Ǵ���s�3I�ΗfEK��Ծ���' �-������f��C-\�Nn`0O5�|���_}d�[f�0�!�f� j��C��Y�����3��z^�lE	8*�R���:�VƴP��$��U�07�Q��H�x���.\���č�I�����õ�$�RhG�����K�7yB���-�N�_��z��Y��ev��n@�k�U�d�ʑA��zb	���.� �<��g�A�x���U����܋X�F��u㺻0��$��.��W"d�_:�,1h��~j*��֔)]X�铷 C�.��\+c���4���rj�f��D���Nl���`�n��{��{D�qGA�֕��?�;g��{�+�:?/Å�ؖ��w���O���qڀ�7_)��V�K�abX��;�Q�~�"�^5�l�!��&6��,-$X�]-�}�"�6I_炟�_��M�yռg,e���dU�l�¡�&��v����C�*�J?�����,��LT��	���~�����Fe"���$W��֕}�OB��~�<�ꄃ\N�n��LV�u-la"�z$/����9����j�9RD�!b�D�w���K0<;��jCء��(�X��fy� ����qw�������1�ْ�'kjR��ׯ�a
\��m�q��T��s