-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
YtxDgbt3m53sFg5LnhhIzxo5UPkHOynbh6BFyYY53lQzT8BFFdv6f/AabUCPTwjQ/0WSlZ3Ewg3d
rRDB6n17+8gV7VBjtkJZycl5N4DBqP7BJzjizogmD+enF5aSBIL/EbyGObQ0jUTMCd68OWiSiRpf
PMHf1oILDx2JzXmOu5v055fC0tkcl1KU1s917tOkQo2x+R8qEcuLoyMXF850jX2uDcOpJp1GTbyy
YEANtLa+hTCY17UXnw/IeBhKeNbSCAiiaIvTRHLd/ngZsk8mrQtUFOegON/2FPxJnjuEf3DluTVC
T80MQElQ4UaBdWJ8LYOQHKtFbLaM/tVabY9/+Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6576)
`protect data_block
dB4gSP1G1EWzEeCM+03g2XaXoE9skvZcFBGxZMftrPqLMDE5qxWh13TamGFEcEStICCdgnpHohFz
woBObRq3TrtMkwscN+daJAR6PMm7eV4KbVMbgxt/zF6SuetCu5bGxFXM85Vpn0TChzUll3bS5LjD
IfAH/xwFWiAXkjLETVJZlWeNjawN9TONVToVUQaAHrYjBBMMQomrwbSIqTNnwXaL0BWlzhCO5MVt
L3VSmhwL0kFPd7Rv7gztlhXxRpvit/VREN9XBLVXJIRH5KQwi5TZwTo1uPB4siQ74hEprgY7hnuC
SwJaJ/tealHM2sr/jIlNviGXIQpztXsygi5g25is5Y9h1dzEO0svp06A7/gvQaR17FHeOujmtQlL
DMHLnE9Eu25/gFfsKZNpflCxL3wJaDgxHTKBVCqGFt//KSOQ8XQeLAGqZ5wD+zSLgTBLL7z4zyzw
vA4/WUSO0oJR+KPsna1U93gUSGItHFHZ5rab8tFBdlsT9cabn3AhUI8G9+0GU67qX4SmrLxngTlL
3feZlzI9kZGx1QcBzMg5nNpcH6Hy2FEpxt4c19ev9YpQJc63Hqc3GESgQXF7CnxiCRht9Fjg49AH
t4Ko5IMzgq6j5gTlbFA3EUl8JEb4lzkX869SagDG8ZyoFZPKazgtAGUwf7HgMXPx0t1drLvvcNd7
9QI4G7j3C2q7U3Mo3EtFBGoh8fBB0nYmp94aG1RJUzpDk4YkVGuXKhc8jJNx0rR/mFJrz22lHDXI
A+OXw1XGBxMTL76DrkBnbtCKjOmJLwF9cDjKkbsX9LxoYSSXzOX4UfWMyBSAxufXSvTjLtgzoYGa
pgHzZOjA051sOoh7qkCLZBmlwIlL8mzVtEPMW7siS5UqDqGw5KYv3+l1ner+7WKshTFSDSF49K84
h3mYi/E5hNhFYHc3PaI3lbjIEJKnUhKf2yP4MgmCEC1JmTlSzysv4vj1vKHg821aqiNsHjh1cBbu
pl7V71Nl3li/VHYGqJJqD2pm0NwlvbPZ4WKYy6pWR8Wf1AWKK5GcqwH/AtfzJqttCptf1diCl0iK
hMdTK3YuB4mdBFGgi+3juB50tocse0ifGK0H3y/W41hoVtAamBG3YhvAgoaU3rOXrn2FmypAPjy/
ICeEAfUF8n06ITM9Zj61Ou7Cv37xhzcIeYvskclQTKgVDqCB0/R8gwu48PZelcHxMMe6/FhzsiTn
AP5l8R9fKkQ4pbkV7O+i/jlIEGd81GpVeGIQ0amdK5vXklI2YuDL1vPueTpFFRfXlzkJVKP+MNzr
xUlPVqxyHY0yA9Pz2uTbbxYEkSair8CBAMHYozsRT0Z54zhmG7BuGgVsb+O2Urw7sqy0ObObc3Vr
ivcZR4TaQ1pF4f3+yTwYG3fOMKi/RH9Dhz7Psi2sRG3VZA+b22CNMCiDA3Dn92SKtpaBedG7AlFf
KvIZGRDCEEu9ZHinbeGa4BJwLvZJPMrFpsDrbNHyHaVbRmVhMCm6iNI0mZRw2ioc7prwCMeecM5P
eGinqqKlfMXPx8W8wZj1KXtcHJYQArWoGEVex5qGrjHj3/2NOpAKMZcvLi0anRtZWZcPmfD6YReF
qY0gzEePZMQdnCjaDQXhjYY+MNrmk74rqqDJIItgztfAQp+ntzijMmtXPsutdSkJZz7Gj48D3oj0
Dn41GooFKcukEOfmG7vHTC4l6ytyOl86Pmtzc6K08IecbCGllheLF8Q1ihLeLmGwfHXXEAcKQG1k
8e8r07MfgThQ5ICY0jxok5V+5UV7PmsRlCno5U3TWZO4XejbKM7/Heg9gXBad0M/dTPqV0Dw9tfC
+UvErf2WUh9uwHHSqfIXLTnGZCP7ehR2LPv/w5UyjzkElu4K8MX6tbLjf75TONM8bniPMznWsFX1
RHO69LNDWz/M1Smn2k5uixeQvQ+ePPMWGgTg6w/XUDCUYfV5CnL/p12tM1uCSt4xaYkdR6iAosGQ
Ss8glShH18BFMGNUmyC59N7fAV6Y+vi6sd4TervXIwHs/BrOnTTNQ/kevLkKO7yfZNlu1WERh5Pt
FxCZbpXZgER9nD6MChKGMcm5if0xXrqZ9qNOB2ll1aLBtHsT3jwmk/B8d1Tvpk7RrqfsbO6mTWRv
TYPK9Ff3KEsMHFC37MgXt0F/ZK2RSCt4GPy1rn98k6R7asG8PcFtvuaJtuXEWn59Plm8k8BNZ07E
SRv9XnZGG/q5k+DLx41DiWzj7HCgh704usC0SV49OvN2lEwshFVakLLUI7KqI2foCfEc7nSu51BV
JwAwjYF5eCWXRx5EY+uNogJN5pfpIznslUHKaXQBNlycX4pk9ns7mEcbE3dS6CLUDpO4m13nTTnf
s4wUMOvjdHPcQluPmWOLTdjGSMcmvMzLVQMmdcLTFr2YeRDa15e474lh74V13Xo+JvARWo2HrhB+
9XLxsTL6ErzHYd4vcDAv0uJ/u/iaZQ/azIKHm2MrSHzuI/DGMxNwIQGv3dzxoLp7kiOnZVoC310L
987PieZhfBgZSjZQHJRa+m0EgQXzZIlM5mw7AxvS4VFjX7hdEqTt1mGRl7n0SnF39+VpDyo3sSjJ
smG7kbMyoXNE+GFF1TJRg85mGEsXewN9mBuk/XDHHwdMOsoZg88J38dSbp/7VE0qhC5vSsnc+CpQ
CQUFOjCK/TJjZ6EuL7z8u8QudsofdZsuVR7JhvI5Ie1lIT0w+SkV811ADRjUjD8UEWO4dsj3KGis
3yj5Oafg3rNpXYPDUbJmxCrayc05Moa5A9Kik08O7EXwGLCm+Jrk3VofN7sSwNaGGN/9y2gQag1t
p1ma2qoq6OTBfH3xR24OsQFXui1WeEaQfKi1KbTEz7V/GbItW89oDlxaALMFgf7fKhl7Y/EgtzxH
/NcUgDBP1jq9llo6WRQkR+1eRt20BJSnhhhxL7VUJFsVJp78sSjzDT6DjZ5DvLccNMp0U7TxDFsl
nTmC9Y+hIJG8XS1BceAkb2OOBtIrWRnLLFwr/9vKsOQSdUyi+A2KGDBcPl4a45tUPS4aeHfEBhdt
unie86sWckl1n0t4vp8JmSzGv3J9VLkBVEzLSEi4rvOy9eXrUBmZlDj5Xr44y7xGU2ZH9wP9wL9M
EuJXmwxkudBy6vHUq/6+loUC7DiKQPRfFf798Q3+bJ46PypGphbWoL3DHJWSqMOIQ68MyxGnhoxM
xo97gzPuFF4NgRCcpfsfnNp5JiJnj7+oqPuXaehOwAGtOnXXnT6vaKFkuJ1wohTnUQbrlrvFu6UL
xL38V/uJdenRiMoBvWSELl193iIoDRGSruFiA6xo0WhKwoKKDZPvM3YEGIDKBVp9NoFhyZoRTiHp
GhvbTXnhUTzT1zhcafGrdRyZfbS4cOT2iz9Cyurum90VYCWQOXqAh9YPJAgIlxoxMOyA3wsLVryg
mwSV6OlDWjTKpmPX2Z/V9hcRDnn5ALCQ1zQPlUlxrpPqxYLl8H7yaZ1RPP0AesnRHRzjEknoEqsa
KTLo4agrie26P8loFQz8tfkstsfmCOyehRW9gTj3bgl0pVEATYz8DTNcmVhRkvNkCyniwRcccBVe
K4kwmEyS5AZQ4ATZxZYQXnwX1A8OhNhpT0a9RUJh8lyFeSbidEJZ9Wx1lkQs47E2DqRQKPu1dSDF
9qMV9OuRtdMegdgi5Lo827VKKB3ybC7BEOXlAOsUmmtCCsvW0Tgk1V3/7wiZs85YDkXH+pBnTuVi
2Ixws5D+WWYw3BRHv2/wmTJjKA5OravqHfT+QZjmg50yC1axJ+hROr/SKodvJR8Jvv1jvgUS/M6o
qvraftHRA13T2iTe/n/jwlwmUYrSdjHp4kghFjk65BULedYGYvVjWRArVRyc+mlN1XVmWDgnTZf6
x8b0Gs26pmRMfbi+NaSgLRwP1eAL17XMZ5GdSBRQppILIZ153+IjSMLIlMYp588rODqVf4TfK9Wt
PJiCKIZDdNTTh0rlEaX8JX3rhYl/Frf/0n7xrODu74SlctLdRxnPAeGiHVH6yQtj2k2Mlmg/bEnh
aHiagMUmHWhGH6vTDBcj+Qpyt+QcN6F2QfhVd9r85AlnpxaF7g3f8eBm+sVRZjW4jsR9irmE1iIJ
+XjetcT4ssov1FR/CzOW3fs/p2P8x0qWQnzaK2eHPBThROODJWIZsKWne+KhEDlW9nrTtgbWBtBj
G7bhdrKlC1sbDiiOm4mrNO32oaljt2jbFp0XCLHVw4/411SUwVKOqz333NOZyhhzeJzP9ViOU7sa
i1FZxLMA/mlyxypIMB0Ugh8HJU07QTpOD7vvSAaYY05utDKZpSs7qVgiKfi2ePSbxJBOnlIR6+UC
skrSZkp7NTJQxVsG+vyM7s72gcXQBCiHQaI7KqZ4o4qhDVJfVdKacBJuBYCtHq/voX3OLhSleIVi
5rEKUvn64UvNBJRsQuhRjGCdbSWNemrZMk9U+NRt8AH8DgvfuueDpxCzW0By0OVjJ7LWPApmrdWH
RpzzLIPH+QXswf8euBiEHTgtnCxzxGhDCnHDuBwoS41blXklZB8C+cBDwkt6FlwckhXulhWOflBM
lCm1KJH0T85h1xljXGZvJPhfKG8godlyVM+PX1knondNDL2hesQKrCenfb8nnlv38QeoTPYqcaus
Zv0zFl2q0jP8+bIxaUOXdQXRHrYr4GaFJ2t4K7BckOlxt8nhpi1EdMQD4uheEvR8lX56sCUeLEjV
qzVuiW9HSDg+cXln8FBMqVmUsikTwR2yxbExNdwM3LTqmbIAIVX9mGC8qzX7C98/GEi4p9wXyxSf
yiVQG3XpKA7rDbKzwo+3ZjsBPOsvqyjCI7jrKgQ8B6aD0LVvudnY70CbJ7PRbsxmbfBjjsNy+68c
GdSG9CKPeun4ARhIkDE6KOe44efp3OXh7/rrWkrl6YaQUkM4zFF3xXVm44+ZF0c5QfMI4P/nVgH+
6EpHuIjzLECDn8m2tWwJYV7laIO0ou4XxlQ9lalxb1oaEXICfR4JGD80j4cfM7CG0AQAgmLq/IST
dshtRkVY54tFHU/Hy//7nbMDBBpDT3oKINLatW8RNJD2MB5JzxQvXrWgapuxCXjrgEjaZUk84Qqm
acHMad0e5I4Ss9afJ2/alBLbyBiHqCmqIXPch/VaEKYBFko/hk0/FO33jHzvJZzqc/tog2kDPTvG
xZpsRhHfjlGyZW9ym/Z4/wRk9IEw/1K1U8HYOGcx1oF19OYPFzLw1MMi2SAW4W6kT8oTsVWjNAlJ
rjTvsdr0JDoN4tIENDyzcJolNDIP1M0+s4WJ9TnvRU52tPUfHU4Y2NsF8zcZwAUDGOqIANhZvTAd
ZZWPs0aKDylaCTmD7n14i09ZJl2BHi1t+H+lVTXdJfN4byfOJfKAibcz5AdFc67RU/mt8uD11jKd
YDxMix91/w/ew8gqc/p9fmjHEg2zKAWio7xEU6NY3AFMCJ0FltI0o0ohJb1iBQyU3CnrDttvKuJr
LX+/wvr2pK50NcDh8Lu4pU/MnIupbGQ08IBK3IYvO260qjoVdVVkR6ogHf0yE8JDAms/IGkfk3Km
gqCxyP+JGHCEMp5PCmWb24BVxeMTbYel2X907/hFJTznzAiLRGrcvmuxu6ZwL5uKZhhlZQFW4c7z
gEOb3vEx1jwbEFzDVdPswImuGlhHZFZ0wM6xuLnsbgMlVnVelZanEsitD8DE542I6Nv6k0y5orVB
YtUL1hP0XO9OPnIGj94d+VWvAK4PQ4Z7DX150UEAnGHnVyHJFnjVlr3f1INK7w4YhUl9ExXK5/ly
U3ORZ02+AEWDbNpkyU+/kC0IYDHhZMU2vX52gVqGRL56Jzen412CkrB3diHkDHl+i8pJoylvcNPD
dPn+6pw+2wpU9Fumbt7MZ4Q+hVQYY1T2j1qRbFnbpCI/erTBi5YLUF+6KSxzujVbsAwqVSkFZXYm
wTB24PBkKKKHyxJOjVMnl09NgV101lqzvmBhP/kjH6krlfxbfqUhkzNxI5uMo0XpNopiqVJpC3hO
Oog0HSSIfxRhErIzDzRtpqC55HUGF0bSAzxxPq24hMwG1Dt9xfgue3YJfbKLT6BviHiiuXReUgnc
IgGUm6aEPeWHiouXzmBOJ3h5v8cim68dyoNT+bxXhSx+/0uek1rU2aCVS7I4nqMp+kY4xdO1u5CD
4wEORAwkR/RADvgK3+26oO+TMo3cdhbA2es11peVSRAmqrjWqHS9SzirZSN0t95LW7Uvk2KzMnti
3Q/U7rrfy24wWTnb84uRjQzD6XDh8DqN106OP6VIP5xKNs7buefn2bEzw1Bqr7wBUytijIeVcPUw
O/GkzZ8t44upT22F0poL/OxL/HmU3QDTlroOYLvEDIhYO3ZOy/mVyemNPMlF20b67P5hDVd3lTIw
/K/0vAxpqp3F8zO57hK9xODRmG7a4EwGUq4enVmvaQgL/aFziI/KTbyr5oqoUvWra8XQNjIWfx+3
/RwcqaMsvPL7UiUcQFN+YvdP0r5rXXa3C9LmKltAobAWUCOTsLIaAX4WN+0UJJou1HW5NgI4B2Ja
592RfqMcODFv2MSMHXnWbmVDrvN69IHk1GSieMe9NOBBKMnarBrybVSGdoZ+eJZpMA6rmm2k61wN
oq3U64pfWFFt4fGCKQa6mcRbbfnlaXFXOolnvuaIGBFHQGoqRc2Y/lzxBxd8vsobDg4nwOX4BE9E
T/0UyoTaY2yVrKWDPikP52NvBf5Zkk2s73tcG09CBySeRgWzajVVlTMWQfKtYnTlAqyggg3xGj/1
dZBFOdDoBz/e7zEC2DQ3FXAlLaMFndE6sPjI9m6w5mpHcs3WONgAC0+pe7cXNfZiVAS9vHDTyzYg
pwtFHQUfFlFOohDjL1YYMaQUGKISX9r3e4P7htdmWEu9CzbDRwLsgn5Ygjr5pETD75Bm6FoPPWXB
svrar3it/aI+2FmTQM8Hv1dCbDk8+XjfIzVX541oYYBjV16hAwTq33P+LEuzAKBrr+xGM9ElOSw3
Fl6bW5VFNfyjdUx2gZFKlLoc+AF3p7uNMdXnTaq/7zcplkazbRtJnQS4aoBHpg9P7iB2YxIKQEN9
tQvfeNefmtokTQq8kvWJlBr7MrIb6nvMFl/6RVZA/Qm9/t9sl3m/662U+cgjTSVzUj9RTfCUOrUU
Pb0DUbZ9f1ryykSeCuuUhR76+ytQgbbQfb6yn8fVYKMK0Ee7puhgBwqHJCeieeuQGfGo8gGyuiyp
LvT1TiIPA08szrRWxvp/edteKbos1nXj9sxzkPC0bn4LXeo6cD5XnfJBWr6M4cKRKuTMw6OkG6o0
j4oK8zHz0b0lL9BrG8ZWyDKRjumpGO0SxFNNr+XlHMFBgcS8SVKDeurYcyQ1wNBMhHibxUGMHI0Y
Rsg+0SfyK8Rsp56KrKP6S6s0LsprvGUidT8y9YVvn57RYLb4teb8MbAz9+tka/+1FEg5cJYIgGRn
hDBryZhL5EBgcvylR7lu4xSYkoBt6Fxn1fR27sn7u1SbrXRkCmysvBVxILgUFRsvK3abjhIj4W5f
0eOZm5qpxpURc2Z9khPzpYxdyLnf3NuoMbDNCkDv/tinjXxetd6hoeSf1bNXsM3xqb1SiHddNO+z
dz5ylqJNrHbPAMe4nJJDsyq0vOmQ6X8RyhoIP7ook+GvKj5KsrM9pYp3VuMU1D56ZRGQjyA5rx/4
bBMELNlrXH7PBSYbhlgJq8QgLCxy2ZIzheNAXVmE3eHftXdEIXwxh83VjGvqUhy4+qFVV8ClE61c
dN2b4ZFjQ0dsrv7IJWaX+sByhTDBpSUJlheB0A6SKW7xRKuNbOGKTAfo6Q+rc11Gim59R0Q3yj5U
jk5viLgI3x4Zyezzy6imeqJKyrMPgQrG22Y36bnIpqWBwfFmRhlfncKhEOkQ2luaeoW0EvL29M76
DrITnz7iym1aO1u5zVA7tUaxoWt/nzZCPHMXpWfh5jkNgiLKLL6ZhvG0oGoBzLNjoOgJJ97x7toF
NNngXV2dlFDwbYkkrg1/nS2w5WIlQ/AqXVegSJc4mxfTqf8L9Q+3/nW15b1zapPTQvxnERa+frPD
MD+ntx8dCGqy+KNK10uc87mzrMsVSdM4KH8TXHdSViXsbGfdI1sgJrv76ICp+z8ifYqfDpkBt/QB
PKAWKFyvBZesc4quwQPwEirFOAcKhWypT99X5sP/uOOmDtkTTHggptUt4Ha8VwGTQ8yDxkHgdMHn
VCqXzeFSBge0bQb7KGECBc6TFOKvuYIlxGjzESyo9k6fUBuvG/UHORca7etLXfgPu65sGTJ++EEm
2ePoPIzsDWZCJkraDZPAWzTABRP5l0ggClUCpecV3wD08zy/3SoslJ/rEy9TFdQAMhmabmPEr9n2
7kkDoHa9Ir47KbP9REHgK2/x1fIZw20zCQDOzInWKdBrlxwnQYLT2gnyXAKOW4W4aiGXgDHqWZ0u
NxFQESI+tJ+Qtw/J+fEsl1es7tNFFb2yZydM2AGRsDIPPJ1CsaYRKC+oM/rswidXnKL990mxtiZU
yJv6CC9ERyki4f6PH2gHtgbMMsChSqR9yI6uJm5hxY3LIwXwPLDAuaimESMfsm4Q2GwMVysu8S1l
Syz8uVaU7uuz7aLzOfcpJWgrmdeYgGz6TpK+rtSJhYGWVN1mQtGy8VB1N4QuC/qyfAxmSZuY8zY+
YrFAhpc90NnSOWXu1Fd6nuRe1dJq9aNt7Jvv14xMaSHYviJg7gfV+thnZXtlxWex7Xy2tAF7EKBk
lP8D67awZkRy95RrjW1MwzQP5ocA
`protect end_protected
