`timescale 1ns/100ps

module tb_proyecto1_parte1 ();
	reg [15:0] a;
	reg [15:0] b;
	reg control;
	wire [15:0] result;
	wire overflow;
	
	sumador_16bits U0 (.a(a),.b(b),.control(control),.result(result),.overflow(overflow));
	

initial begin
  		a=0;
		b=0;
		control=0;
		
		#3000  a=16'h2222;
		       b=16'h4444;
		       control=1;
				 
		#3000 a=16'hFFFF;
		      b=16'hFFFF;
		       control=1;
				 
		#3000 a=16'hFFFF;
		       b=16'hFFFF;
		       control=0;
				 				 
		#3000 a=16'h2222;
		       b=16'h4444;
		       control=0;

		#3000 a=16'h4444;
		      b=16'h2222;
		      control=0;
		#10000;
		       
		      $finish;
		      
	end
		
endmodule
