��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,<�#�7�mh�NB80�0��Q��]�N��5������N!6:x�q�!8�<*�5�)dk�r?���F�|IY���IА]���^��h&�V�{��C6���'4R��'�yd��r�����ց��i�G��9�	7v`53:��0����a2��5�4e�T�˛�����}0�+��e���=ۙ�����.(����	��Ѐ}g�[�Zv���'XЇR�����[�:�/n���%/��&˵�(�Aa��m�l6W.�@��D�t��:�o
,��x����E�������ˍI2)�x��a&;W?"�+^�X�4r�b�I��~��W�}��d���}p��y��ٓ�?�z^�5��Ð���*-Z��e)��t�9r�>�*���D������__�n�E���8 j�+��WaD;Qc�"�u�~WJI������'ʖ �<�=
ڈ��.
�nIS��>�P"=��R��g�Gͷa�59�x�W�$&,�D���y�� ;�b�v�� �Wh������Eg[� -J`��8Y�Dڄ>������[����t�U�{�PB60��T n�Z\��O�M��ӻ��0#�$)F��C��k��w$���e��m�M�ӞY�GcS�~�ߩ<�b�����/�u��l�z��4^��Ppm�ajIP�=s�{�s�Jp>yvƖ/�B�_��dx��.����*�#��U�h)�c����jg"�)�r���-U�D��sKT^:ο�\�1�ϞU�U'�CR /���r�)�Q�%�� ��S��ů����5H�r4{0�vͧ��#EH/��#h��Th�)�zr�s%�$$�����>P�