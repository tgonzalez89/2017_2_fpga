��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,h���~�G��G�j�V,=�ԸL7���[��"���:mL�Nn6?��.Vts��$U�S�C��I�i�j�붃�}즊�üå%����6W�	����:�-�=>:s����u
�I��3�G��U��Q�����I��F���bHiM�x7�$c9�ת�cI��h���5rTTg-�z��;5�CkB��f��zI>�p�8D#���@29�h�x���{����r����`���\-������)b�-��g��O�T
$q���R��o��H(D�S�q�����:[�px�b�� c�`=�q��k���,!Ush�o!��4n��j$={P@.��(��\%p7���WA([�y����w����G�_�I�'���bw�|��v,Qm|0�I��\?b�R$ײd?o��d7]h�!������O=�Bd�U��>�Ƿ�H�en��j��6��鄂��/&x��A+�P���WJ��+3�"FV�$���m���E�T�%HZ,���!��3��Ö��e0Pm�+!s�p6BYx�z���E^lbu`�)Q]��B�@ju����;��9[�p����l�b�x@�8��5����VV��@_��M�t�H�Y>�u𥄻`�a�q V���4���mf����VM$מ�B������O4M� �'ի�'�?���Ì��9�������R�f6��q (%-���*R���d@�Ql�2:���Ì(Sr�pbS�n��e�u�%ں�{�I��,�}�(R�m�2����R!j�w�
����/����_G�	�_m�0�m�� �5L_D�������F���i�>�[��ҏ�BM︡��%�`?J�G�h�`�B�6F
�
c�OF��?B���]��K�\,��f��}?rE�E`�y e��q!��,�@r\�a�G�#uR�t(^�H<���E�:n�ȴЄ�A\.^��{�J�ìRoSa�����ߞ�&���]En�gY"7��4*���i@j7�i����aZhoB!��P�����o��fl�&I@tz	�ERk��-�(U�֡'�������\lѥ�����"��� ����W��V�;!I^��L
?5��P�.��� gzh���� ti*�WD���	yaISn�?[�h[xG���Z޴���B��-]Wi�B���@纱z�K>H8Ⱥ�Z |�2���Wd 䗥��4���.�(�uo&�52��hzw�S�����'hc,D*��l�}C�Oq�2+��BFp�=�ú�\������ި���A�U���jVL�����L�����N�{0DלN�J���|+�o����B����s�s���"j*?�z#�Ƴ�xc�ɣ�M>��M��1�d�F?���X�#�wI���D��#5/�;��A�����0��$�@:	TI?��@D���z�r��Q�:M��F���g�XC���>�����V��l� B���v��YT��q0�2wo���z�x��s��}�G��3&	�x]�!	$
d�_���X���R��Ĥgc�ii1y�"�NSv۫�JDu���F"<8t��Ɓ�yW������!U0!��V��Q���b9??��CH�4[����٣����R�b0X�>� �q�"t5��u�ȝＺb,p8���@Z:���c�N�;ZR�D��w�6��O���:q��n�2 M��)��)������Y1��7#��`}�	|�S[�{����a�Ѡ@(�b0ݹ�Ask���^I�W�R��O�hg��3x��ҽ��`S;/��u��;̞}��^.�Pw#��r�iP�T\7p+��ـ�Nx���Yj�
".�!�r�a�4q����S�������>@"� �I-��oZ!G�eP�| ���gw��X�c����w��o�߬�ƿ�X�e��hֈ�b��G�l�&�u:�\�w�Y�'+[!O�F��Y�5V���氿�$Ā���L��+���K"$����45q3���r��T�DQѯ�\&CKߟ)=t�<���p8����F|5��!g��4b{0ɱr՗3�`M�����9��f�4��~����=��'t���Z Ig=�z!�o{0~�3���ᝍVϗ�/�\�N����Vm@��	�n�1��[��f����c�۪VB��x}�ԟ�{�~�]��M�5��� ��5�hC*���ᦨD�Zĺ#���'��<`�~P��FѰy�?N�v=���#��IV����]b��R���ԋ�K�5���OW�5�U��>���
/hV�KH7X2��k-�����ژ�q�nV��[�<��}J���/l�XM��1� ��"��	|�xټ<4�y�#M�3�,,�g����>^F�;>]u�uSRv+-�	_4�B����0��������ݺ�ֵ=���j��iK�1��B溃=E&��g�`�6yN����6���#���0�+hp��W���rd������8�[���:"� ����Gp�l۵��j��5',X��8��ŬN�����+��>��~-lK��������	�`��|��!�b���>Ah���x<�M�.��aK��
���|z�o=
B������3/�m�駻�5��֟@��ފ�;�H�Z���/"Z�B�㑛�o��'߮��)��
l��l@��b�o���Y���_j����wS0�(L����d��V���'�-�E��y��:������x�����2�������^��>��(�T��h���U��'�TH��I��"�٦�J�.U=�[���{�{>M�i
����QN<�VjI�(Y�>�+@�J�d�aIW��u��K�mtPԗe�ި*;!��'i
Pƛlys�����uD#�:��\35]�쐚�t�,��=z#q�,��ڳA%���p�{,��(.
3�<��w���Mu!)�2����,ŴE&�U�U��YCQ�Lf	n%(,/!��������7������� �(p��	r3��)���ߝ�b��	��8�w��NƮZ�<N�M"� ��~���*�Y�/��n݅�tˡ�#�E�R�eߛfɍ?g��Q�#���)�m0X��
8�I�>]d����k�Q|r7��s��xy�T�q�m}��/�@�i5E�/��k{t5�0X���UG�%�OM�}��ԧ���]�'��Plmh|�U���A��8|� �Q�5���P;���du��-�ҽm���9۰3|�F�qr��+������E#XdNS���G�m;�]1��p�$"B`E�!�ǅ D��yC�� |Y�|L��8��J7�s���蠦jy��@y�p[��<%F���S�z��b��A6���#/1���ݦ�u���hXP_�Ǥ���o$���
������N�rA6$�Ġ!H�3�;M��r�o��.��{p16�Wms=�ǹ�D!`/*Z0?9���_
�f5�
�O��J�L>�U%,$%~tS��e����OOS�F�l�)�~vz�)+:�s��}.����=H,U����KqBT��{�$�Cu�M�/Ē6K�$X�<��w�/zƪ'��O��컏j�!,����r`[�8��G@�����P/�~��C����B���U:��28]�\�g�Z���_^�6)>|�[@�EK4,̵���z_w�����ZA�.�g?
���Pp�>oE݈�Y�-������X�2ʟ �k�����)��#ݾ�ϸ�Ab�f���+�&���Il�KFw���]���o�� ��s��i<{����9R�C���;�-��՞��%�A�"��<�*�vF}�[w�	�M)���d�i6-&�m�#_����o�@�<��i��ýs-�L$���r��yIc�r-5�dtH� y0���SN�5|>e4� k�.�i����>�|IiQ�f*.oa�U�g�n��Bi���E�):�B�4�#�vM%����hpM�;��w4`�}��^�R�4I�6��%�y�j�	M?L���j��p��ٍ>�Oi��گ��*�=.}�,i���wǈ6��'�]P&�[xp�����'��#�$����$�ԓWҘ���O5B;0mg%iXdӌ#�5%(D읾,i�a��5/gO\��^uzb����+��O�鼬��?� �����])GTQ�P���h�h;9�B������_��.�����J=����B��������%��U�sx��p����M�+�[γɩ�������,wU�XwU7a��������w��j�nl`�[���̒�q���q%u�or�:�tl� ������]89f< W��V���f���a`C"��l��S �]�g�q\J-����-:jH�aGv�>�H�����d�D;�5�J�`�6U�ܝ���q$(n�ɍ=�M�����n���f�݅��w�6�Y?��D��%�ȷ󑟭Lꂤ/���R��&��47g���f�]ճ0�k�,�8I�x�gө%r�V�u}a��mX�Q�����$-N�P��L�[��VĠw%�5Ơ�~�<��7���9�}{��\.uYY7Is������c'ez�7��R~��p��Z��紀!r�Q@��9-�.��������~w�8�]4�r��+� 
d���*�3�o�b�t��s�J��mU*Sp�6�@���hJw���B\y��`v���������#�fć-�/��K�\M�/O�9z�����!@YU�6�:����x�u'�_]�zt�A��+)_G�"��y��c7?$�ƋG��m��ś̨|?\�E��F�~�|N�+��Ӱ��3�	i����I����Z�o\s�+�,ځ�_./�� ��� �v�������?�|����K5��!��%�G �'<�J������_H���#��6�0�����
r�sܮ��j�Q{���n��ˈ�&�n�-E�ZN-$w���������S^��_ZN\�����#9�xh����W�������RP6	�`���M���N��
5��N�+5�PO���Oo����G����.&�`��!�Ln��x����c1VB�/?u]X+�� ��f̾��r~����gw�42�,�)q�T��c]%�m:N��c3v