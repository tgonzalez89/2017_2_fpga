-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
LwlibNCtfhb2rLYkKgPVV7VLH1RXE+bd841rqZHWWSkUfPxP4se1Ef4RylkNFk9jh2HCR2DkVcT7
zgU7e6z6KODd/Qa7bDTb9X5w6gifbXGQCpG2Bak2NqB3VqpFlKJJnXQ/VFlSHG/3A0arhhVf4h40
zNC4GRLldNh2JjLGANz81w4V3SFMMvqpWG/N/PfjSYkIM4hba8+owKxxbYu2vLnwy150jjLN/cxT
nhe4wVN/PioDY0H2EI9n2CCWjfvSvCBpILznZvxgDnA0mO5zGpP0mZSgrOrE2dvV0wHMQGbzfqHC
8lKXf2PJwcIlwMfrFaIgCEPY18AqCHxsX8uxQg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5392)
`protect data_block
uzgA+j4ShRaUlz/Z2nZZQT7mt/HzI8ICKaW58o5ZnVN3eWql6tP5uN9m7sY5gFi/eQMlOHyeIC1i
rq3bEQHZU54tAPynlWOw9SmGATPVjq/ipT+/PBgXofCSCAp6gc6jKNxdnjMHftHl/mqoKje24bO0
s0wpjm0A6Sl8JW5uBdOK7gMFYv1TckByUoqhDkohl9HFuGrGwS7ZIKVvnbwv6d6O/vUB48iwa71e
KgSbeXT3sgu4HLBS7Njcwj3u1iEGR1KB/ETFbVTHmMJM+/MGcpNReAXhf44jimNC7q3xPrOD7I4a
F6NByHLvz0QnSU8sdPQpezcNDDNqdSj7c1dRQJIxBRP2Gyv5jQ8Fp82/1eXxTzO6GXZUS6Y9C19G
1eweBq4Nmby2fvxFj7MUm4tlUFwMT6tC7QyvI7jQA7jLyeNh5WQku5wW/8SImpJz5vEYyLelLkpj
BqaeR9e7NTQgKklfWZTHqOQLjE0rQfzHCfbw9oB3KPVlyRoj3619yHAdSwCGhyGAlFLbzt/ObXMA
wbPfvzGlsIlM2DKxww5r5QoTuCZRKtUNjlIwY7FmJp426yJU3ylExkIceSI0S21fFYcQya00NG87
HUMbMRBuglYLC7QkTYqcJTAt0L+//LaxaSxZEO/1Tq7gtkEULvwBSq29W/Q6qYfMc1NEnWmODNKI
B37udxVac7/l21hWNyWy71pOX3dP5KcYCeKte0qFFeT05nkk/RwfaU0maO+ULeSJ8wNefuCXNpUh
Hs+aqPGoMqIoP3rYBuRX62DMNeZ5HTUz4RNemYXXoFsEV2iFBNwG+N2et5ztvQWYS1pKe/fJD3nj
nrfF7t/F/3aqiuUcBSV689yN6xiKMAi0dPPCiHAYugMG++Nqf3zUAhkr68mIDnCCz92tp7mqP8Df
hyLAydzBd14Dw9VPCddpw8jmZTOXq/eXIpgEJmb0tIE5AK9zEpeqCHWPZ+UAuv870x8795gPaNh0
lraTRMaJaAecJbTHPPVJaO+W4MySq47vPN/ZQ5eZnPgt7rNwTvAnKeMD4q7QMIRTC+7uQ+8XN4QG
jQqfX7Az/s3xSL1HWt5P6uHQ5228vrf5m95STCmYFqEQ/dmjpUg8VS2Xy3RhULckZBAqPPeSvIVL
DoOLXds4hRJoXvPKh8PBXeRH6q9z97jndEQBKbv7iVQ/AVPPHb+VqoVUShM3nUvQ9CqKFMtkUvi5
DI5DoLJYdMVoobuO3CHpDdks7LiMqUdBkAKqbd1bd1QQ1UUXjJZdyxUGfsufDfjzX2vHiuD2Mimq
OvH6QTYzNxOGgm2XsB4mcMwaxsBTdNfnalshTuG61rHJd4UTWpPkYoYKqvSXPg4jspJFkkrcmNfL
UQn8gMFGfmrw5hd7GJBQ+fwuXAIciQqWxQR5I1p3lMb/pbcpwRbZJ0Vxki67IF69OfFkvk9ll4Jn
bFu4CLG56AFnEHMxdU8OmXseR03YWuupzgTza1biHiP7Sl2eXzteDlkk0+SvNsB2wB1fsP8i9Zpe
QNHBNFPh/zEPB9gB5dm7y5i9UYf8/zSrF0EBlXrrO7GiB2RvKCWJh1pvl5ulfdKT0StSclU8v1/W
i1DiLlEkDfP/QLoUzes366QsOgXcF+/QPq8C0igmJq+umHmJuopkwrhouunugBLpZmQuSM6EgODN
Akx76ZsFvSR/jfrhXI+f3myo+tPK+6UrwUj6waX3G0bW92t1zHFLZZAc1hplrW3eNBGZBC5t1q1J
19XyebCSUGD2X9CLIi8zj1rWQof/ngixOihvBQNybSEDiTjlHhHXlJJJhTceFRxRW22Tjbd0G081
fhhZMBqzNoopLyGZ65RT+b0HwTvQMr43uVSNz6Yzhn/xP3koTEw68d8oRY3pVQyf3udS/6RMnFmA
iCCF2BW93vs0XEjepONS+gkIEsuO5MgMrWZEdA64jyQ3F95dssDgUQqvDr8+4zSEQQJT0AcBr1Gh
/MUFjvAz/zAzGSW2MRH1Xb79Oi7U9l1cu3ppS8Drr+ictquJBBokpv9gJcFl2plwkSpBr1qP+e8Y
J+gzk5RCAlzUX7T6m4S5DVgfFJl6kY5VkrmRxDqR1h9HeV+eZMeb7uLZtdzfygsu1q2kC8k4jGai
D74/nQjTici+jyf87tO6Y0+2BlyB7YkecYbPEiI5HeP+2N2eG3kAwA3dhUinB+ckFHGoWwhv6Ole
Zl1Q/1DPQAG9rv3BZKxLWl8UeVHFB7Ql9EHsPooCcLd1Yvs8zjz7lw/8PTkU4JeAuT8O5Zt8jc9/
VYWR8KqBXZZ9I535qIVowQDgvXFER/ya5bco3kkGpPzwgehuPmANt64OIQG9urO9vXJuSZaoyejT
fglQNcxsCfPNzdPUIUHSrPFlbCQeWQkTu1jzv3eGKM1khWbccynAzH+451H77NuiZ2CTM4L/KhuC
2flJE0wSM4nWtJR+qfVjgL50R4KM/JHThlveaG/YSCP/UraDTiXSS9qWjaN2vU3itPByMSJmonVn
7yVxkONcGTZx905BSkr/BB+rIx029vfVWmqYPuRnxbGXSRR8rhYtwENm6niC/h9Hes1otDHIwKsb
T7xF00ef4oeZD/V2McrdT8jXLF2P+tJyfjkP3xfTkxkr/uRBdYUFVI2f0Va/aEjHPnEUrVmXV88b
+nuy65pMkZzEj5C8wLGIq69ogY2bnc4w+46v1W7Lr5bPCQXbAGY+UeqMIj8fN9V7ZWpyPsy7wemi
LFfLPpQT0XetPbqDcHZC3fsRKU3tDTQSS9vuclSmDZDHDtw8JTY2z0kP+zqHpFimk9cNz1djoFDo
xJHqxJgoe3V6WmmxpLzx92ha3jTJSBUFoocvCKY6YYWethcLQrY4U5aXSzX09m7NkzdoaMo+gIR8
ZJlEzw4UGOGRlk1W/8bVm4rg4plHS5kcfm8ts7JrGj95Ea4cFJKGC57VJUDy/VyON5DstEqmUel4
SiwNQ79S5wx1++zY1JIgoc/UZLRfSKpCnv7dySGXBWAzSueVUBgjQ5bRVMGrheqVJXr88+ejKT7f
awCeTpculAd+i/H6gFBRtpeQq+JTMNnOyzNuZwGrQUatxgmSzBKokZ721SHjLZbvyYL+LL/dJiop
ppgccuo9uQaBn2Mt7XjWm/DubgJjCRurGrF58sx5A2LFXmM24y/0ISzvU8pEZkQx5Hdh8vdExR64
G2uw55bT3uPi8Sw9oeO/GR4qOFReKyG/skfcWtd1dCDXBTSgJStNo/4WIwLtE5UaX8JQDQ3e8Vl/
tq20uWIa7ePAQHHogaPr2b6W6MHaXtiMp+yaXBPXCqPE0Y8Y/pWXnlTuEA4buulyOA0xqmLBJgxw
d+D5kgxfAtg2wrIqREDYDxize71lHwFvqFillPcuasIu+LEmw3V6tfADLBKyNjqVpaEyyAYbOoUw
HeQwzj5c9sV9OAfiFe2wm2e3lVZHfOXQw9GC+lP3GVPTFXMUXdhzfpvJubKUK8x7Ope+6wV1cBnQ
MohTvGNQjkfs6W30yXG9wgF8EOiCJu1Ful5WoDcu/nO1RVeplUc9rQnet0ns1n+uT1/1TRnvcVV9
MXtMIx+LsriTtmO2EP8jVAtVlv1+aBQ04qQ4ndBtX650jkPd3ubvVPiXDh+wFlyrkKSZiciU/kFJ
KYUw9XGVjU0fptckLfg+KTKMP53qRuEj6b+YWGnssmV4LLcqnR/ZffcmIQeCrQeJ9YzNHRGMgskA
6MiG14XhGy8nBCVycQmqSHAPzPZNfGR4zUUGg62CuqvL76P7hcHxs4ow5uu5vAh+0MNWngkXQxQL
EDIAQo8gQg07w8Z2xnwo3sCmkMD20CQbm4y4Qro7F+VtgG/gWUpSdPgfjX9qwyIjFUvztpiMkbTD
eTDqFOmC25yCnfBXE5UMUDifiuvQAaJi562R97cjZN6TOFTVpx7qbzCXqRATAD+dkxofq9ypzeAi
oLBzw7apaWw+vtNgNujr2evVcIdd0mquF/E8opNWDDWGMkHLrHgDJXmF+zeMmUCY36R3UQR5lMAz
Od+fCOdF+vRjNV00Cq+fl80aYhOWEtxM4G1T5wkdyMdAGXZtd00ugUfdiduAjZNtkCJy7cLuMGKo
2hDoCxC/M8nIp/ta4Q4AXAIkrw9CSMArXAr3hiup5/JMMsp+VkywVvCqVfhJ7dM3RhccRqbOrvlY
5NtTck1mG891JVsnyi00wh+SxnkzG/qXTOBzTdrzs71HeytAa23bPm7dXxtFc3GqisiSkgOO3Bo0
8FGEGPJFgOp51s79jO6SWXlxMI1Etg9qObfEGy/LKI3bpfO+BAE3Si+aQ7iS42PwHeULAAMV1byS
wofGemmwTk7CdvnP8ipJNYhdTXnpgdcj9xxOmAKNuSK1B79XvYmh9z2B4G2SkaQYBFBJI07J0oM6
PpQnSOW+aKYkJR8Q4pPsn98qarQqPuf/d5yGTA2FmJFU/g/3gNY9atXJFKWosI0U2B2IbDnmTofF
NSQKw0ExNQyC92Jonq5J3wh/WGpsauQ1pxCQhjs/7piAOtoVp5Mq6g8AfyjGaaDn5dtrcUAwbaDJ
G3kNnC9B5JWoNqWEttuEQ79LBFWUWn/oomIboojCiBlAQIHvme0hZaP+idzo2u0EcJHe+M81nbMQ
mvpWwyeWvaEcYhzpbuPNptVy75MrfS/xseiWJRRsXws0UDCoPH8uFxBz1JRkJ2iLhZ7EQnTKH+qz
mSErzLMyIx7cpggEV+IvIRMA7K0iONDIYUEZMrjpil/fKA2uui1YTEd6NUiI2kIhT45enwYgBJlx
jzpMyeAleftCfxsm+NMIlyqvfc5qktDuIrcdl7zfPidSb9kumVOCHnwpl9t5JgYt3ymxTocrQvul
08LeVD4220In++RjXMr/L12EzYLO6Cef/1JTd61NzMLS+B8fwCXuvxXxPcaTZDHo5H/3vIi2Qa3J
QmQ90FWf3vN2ufApQv3CBuo1O4nnuB/kLdvGkGx5mggPhSB31MzgR5m0JPT87soh6pMy9Z/0CwAy
fp97y9iWAHSCB6rJosWRja0BytPrhEnMuP8Js0P7VNZ1uMDpkaxmQMiHCscmiF23llNI88KhiPfL
dUbrJEA02w183vhyYpuGFD7rKyjl+S0aeKadtDXuE1owByRYF9qPqby4Kc60XekWeS5tpJp2aSXc
3D5t2QgFeH3T/6G+zS78vuwcVG5FyuDCKGdPBnU/r1rqZCoQng0FQmCSuT2Sm9pzcDTgPhPyThZr
SKb6AHSYrkVxeGhPdI1DQqZVplVSDn6eeHeFnm4kdY4NbomrPRtCh1BhaVgMCuUjzGljMYXYUsAl
F3bX8zjrAIXjuBki3x94hvbKemoCq7NdtNWTJTjeWyHaG5GCtBcbGlGi8Jm/Zv+i94Vc80hUwBGr
kH62y5AYDt+SvJk/Vi8F/dDsqVlEaNp00ebpwzTqPfssBi4wglo8YKIP44tnLJA27aN8w4zZFKJd
eX5nM04zzXQ9piGip/SSUMOgh0NXMi2WjKO15uSFEP3Zq8qehq05TcXvKonkcSGVacoDOoCxm8ye
VpPu7zEjREYp5qhHYe5CuJrK2EXosSrBKZOSjXH+58QjNCevKqmniflZUTMtRxXq0VfIBjOrqWSb
C/9e0SnDmYaDVXgb+JJ6/B7r6fYKGrI0eQPwC9XA0W10iTBJOHiSZ0kk0rJy/Pz9JIZS9QY/c2wc
RSlr0R659sGSpniRc2VoHslnDNWEOpdHRmSxtz9qfWkyIcgvnDiyPpS2qINblJH2ZAo2cplXXUzH
pxQs/Cfa7MpzzmJhLyj0ePnHmbCpbjherKjmMz6Nei3XYbDLdYhWV256jejh12oQXQXhWf7E2bSO
Ga6eZRh/HLvnSHKI5r5gfh0A2wKlSnImQyqIsYBVVDo5nU/WsgIx6PfA9cCrOJlnp2V+A4fi4pvr
2m4mrGOz/zb+k1C9/YjADhD7CzMycwrUfeMhrluP/lw+yLXIM5/MYBfVeuFoATrc5Ot+e1whhIPw
HjB0KTzrqlj21f2Tg+1RqzlGjM+89Zm93uOLCNlg2Eyu+gnaK9lwFIEfOqYhQPDr/ijNsx2U6cyA
kuo+oEKPmXVzj0t3oLM/UKN2nMiS8R8pNE8/8qkef71y6b8SkAZcUusVw3jCFbBtogLrv6fQFNF0
GmBp6tukYTQIaLP1Ku3vFiYIg1ub1Fv8sPM+eI4QgjjUo5CWHy/tTPGW0669VzkHjji8zejqjtxv
9neV1P61Lk8o2z5fDNDY0v7D2jHUnY/zbKbyzn3gmsX5l8qXpLmRvjCbL3EzsxrEaQrnayHCUBQH
mJ6jKOJ1JFJ9v0Dg6E05sJ+cuBCeVDxeZk/4mQimRgjpZ+h6Dtm4L/OxnipkrGb63ViGJ6y2V4sa
ODo9O4/KyC8FOhDXUBxWACuZvNKJkKA81d6rBnJm3ILwv+Q76freZAMxS5vf8mvCt6qv0+GXQVbY
c9SqY0Hg47YybQiMqfTwStcRtrI2+wDWvyaXh5op8Esh4+U3rJCvaHyQKhYpIQ4ai886ZU/fcGdp
8MU+ENT/dBR2iSnU+2efBkv2RTRSlRc4nzSD1SA5jFOYTsp1LPy7BZx+M6vplhoOABjKNS/IAD1D
ERYPYjP49YeUmWqowY8dXgRzwDa2lKlCf2uZ3Cbi/eWUCDomB+4lvcMWn4BaHbOTGEsLOERQGXRX
E7gfiP0MoGVgUM7sABz/3fnAOZaT8nA1Ce8myeHiIq20lFekjrr488j9tysT5T4kuf+UBJxvbJRh
1VoAPEL0TSkUQDWBMaRZZEhvmjjJNfTXt42UOjqKyQWZTxHV6ppDqLYKtUGQN2xT1DalZqwapBpC
XZrmub811t0YkbX683eVZMW6cwHWfPhbb9q80c9ebj/QrR99aOTnPL40gn8ajoThXz7yIEHnrtEU
iXaMe7ZOcL/8Mv9PYx/uAif/KInLuSnvfh0rpK5xeNjpdNsutKhMCnkeLuYIFSqLcIRHAEtSgbNH
PaVQxQCWvhurHmZLzn1sTrXmWTmRB+Bixx3yko3ASai7Uj8uXnFbzOYfxGlNEM5xRmR36PZHp/gG
lbYhBAgCyxVAjZvI3QQYQFtkd7xtoKUZVSoF6aC4+orWUdaCAhMq+vdxIY4n+nFOUR7Npeeipf6D
XGc0MuqnK1BzXR2RB80yXGjZbvoHQqZAec/RQlMTS1x/sA==
`protect end_protected
