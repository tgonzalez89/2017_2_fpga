// proyecto3_system.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module proyecto3_system (
		input  wire  clk_clk,       //    clk.clk
		input  wire  reset_reset_n, //  reset.reset_n
		input  wire  spi_io_MISO,   // spi_io.MISO
		output wire  spi_io_MOSI,   //       .MOSI
		output wire  spi_io_SCLK,   //       .SCLK
		output wire  spi_io_SS_n    //       .SS_n
	);

	wire  [31:0] nios_ii_processor_data_master_readdata;                          // mm_interconnect_0:nios_ii_processor_data_master_readdata -> nios_ii_processor:d_readdata
	wire         nios_ii_processor_data_master_waitrequest;                       // mm_interconnect_0:nios_ii_processor_data_master_waitrequest -> nios_ii_processor:d_waitrequest
	wire         nios_ii_processor_data_master_debugaccess;                       // nios_ii_processor:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios_ii_processor_data_master_debugaccess
	wire  [16:0] nios_ii_processor_data_master_address;                           // nios_ii_processor:d_address -> mm_interconnect_0:nios_ii_processor_data_master_address
	wire   [3:0] nios_ii_processor_data_master_byteenable;                        // nios_ii_processor:d_byteenable -> mm_interconnect_0:nios_ii_processor_data_master_byteenable
	wire         nios_ii_processor_data_master_read;                              // nios_ii_processor:d_read -> mm_interconnect_0:nios_ii_processor_data_master_read
	wire         nios_ii_processor_data_master_write;                             // nios_ii_processor:d_write -> mm_interconnect_0:nios_ii_processor_data_master_write
	wire  [31:0] nios_ii_processor_data_master_writedata;                         // nios_ii_processor:d_writedata -> mm_interconnect_0:nios_ii_processor_data_master_writedata
	wire  [31:0] nios_ii_processor_instruction_master_readdata;                   // mm_interconnect_0:nios_ii_processor_instruction_master_readdata -> nios_ii_processor:i_readdata
	wire         nios_ii_processor_instruction_master_waitrequest;                // mm_interconnect_0:nios_ii_processor_instruction_master_waitrequest -> nios_ii_processor:i_waitrequest
	wire  [16:0] nios_ii_processor_instruction_master_address;                    // nios_ii_processor:i_address -> mm_interconnect_0:nios_ii_processor_instruction_master_address
	wire         nios_ii_processor_instruction_master_read;                       // nios_ii_processor:i_read -> mm_interconnect_0:nios_ii_processor_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;          // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;       // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;              // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;             // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_nios_ii_processor_debug_mem_slave_readdata;    // nios_ii_processor:debug_mem_slave_readdata -> mm_interconnect_0:nios_ii_processor_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios_ii_processor_debug_mem_slave_waitrequest; // nios_ii_processor:debug_mem_slave_waitrequest -> mm_interconnect_0:nios_ii_processor_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios_ii_processor_debug_mem_slave_debugaccess; // mm_interconnect_0:nios_ii_processor_debug_mem_slave_debugaccess -> nios_ii_processor:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios_ii_processor_debug_mem_slave_address;     // mm_interconnect_0:nios_ii_processor_debug_mem_slave_address -> nios_ii_processor:debug_mem_slave_address
	wire         mm_interconnect_0_nios_ii_processor_debug_mem_slave_read;        // mm_interconnect_0:nios_ii_processor_debug_mem_slave_read -> nios_ii_processor:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios_ii_processor_debug_mem_slave_byteenable;  // mm_interconnect_0:nios_ii_processor_debug_mem_slave_byteenable -> nios_ii_processor:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios_ii_processor_debug_mem_slave_write;       // mm_interconnect_0:nios_ii_processor_debug_mem_slave_write -> nios_ii_processor:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios_ii_processor_debug_mem_slave_writedata;   // mm_interconnect_0:nios_ii_processor_debug_mem_slave_writedata -> nios_ii_processor:debug_mem_slave_writedata
	wire         mm_interconnect_0_on_chip_memory_s1_chipselect;                  // mm_interconnect_0:on_chip_memory_s1_chipselect -> on_chip_memory:chipselect
	wire  [31:0] mm_interconnect_0_on_chip_memory_s1_readdata;                    // on_chip_memory:readdata -> mm_interconnect_0:on_chip_memory_s1_readdata
	wire  [13:0] mm_interconnect_0_on_chip_memory_s1_address;                     // mm_interconnect_0:on_chip_memory_s1_address -> on_chip_memory:address
	wire   [3:0] mm_interconnect_0_on_chip_memory_s1_byteenable;                  // mm_interconnect_0:on_chip_memory_s1_byteenable -> on_chip_memory:byteenable
	wire         mm_interconnect_0_on_chip_memory_s1_write;                       // mm_interconnect_0:on_chip_memory_s1_write -> on_chip_memory:write
	wire  [31:0] mm_interconnect_0_on_chip_memory_s1_writedata;                   // mm_interconnect_0:on_chip_memory_s1_writedata -> on_chip_memory:writedata
	wire         mm_interconnect_0_on_chip_memory_s1_clken;                       // mm_interconnect_0:on_chip_memory_s1_clken -> on_chip_memory:clken
	wire         mm_interconnect_0_timer_s1_chipselect;                           // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                             // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                              // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                                // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                            // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_0_spi_spi_control_port_chipselect;               // mm_interconnect_0:spi_spi_control_port_chipselect -> spi:spi_select
	wire  [15:0] mm_interconnect_0_spi_spi_control_port_readdata;                 // spi:data_to_cpu -> mm_interconnect_0:spi_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_spi_spi_control_port_address;                  // mm_interconnect_0:spi_spi_control_port_address -> spi:mem_addr
	wire         mm_interconnect_0_spi_spi_control_port_read;                     // mm_interconnect_0:spi_spi_control_port_read -> spi:read_n
	wire         mm_interconnect_0_spi_spi_control_port_write;                    // mm_interconnect_0:spi_spi_control_port_write -> spi:write_n
	wire  [15:0] mm_interconnect_0_spi_spi_control_port_writedata;                // mm_interconnect_0:spi_spi_control_port_writedata -> spi:data_from_cpu
	wire         irq_mapper_receiver0_irq;                                        // timer:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                        // spi:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                        // jtag_uart:av_irq -> irq_mapper:receiver2_irq
	wire  [31:0] nios_ii_processor_irq_irq;                                       // irq_mapper:sender_irq -> nios_ii_processor:irq
	wire         rst_controller_reset_out_reset;                                  // rst_controller:reset_out -> [irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:nios_ii_processor_reset_reset_bridge_in_reset_reset, nios_ii_processor:reset_n, on_chip_memory:reset, rst_translator:in_reset, spi:reset_n, timer:reset_n]
	wire         rst_controller_reset_out_reset_req;                              // rst_controller:reset_req -> [nios_ii_processor:reset_req, on_chip_memory:reset_req, rst_translator:reset_req_in]

	proyecto3_system_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                                   //               irq.irq
	);

	proyecto3_system_nios_ii_processor nios_ii_processor (
		.clk                                 (clk_clk),                                                         //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                                 //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                              //                          .reset_req
		.d_address                           (nios_ii_processor_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios_ii_processor_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios_ii_processor_data_master_read),                              //                          .read
		.d_readdata                          (nios_ii_processor_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios_ii_processor_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios_ii_processor_data_master_write),                             //                          .write
		.d_writedata                         (nios_ii_processor_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios_ii_processor_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios_ii_processor_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios_ii_processor_instruction_master_read),                       //                          .read
		.i_readdata                          (nios_ii_processor_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios_ii_processor_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios_ii_processor_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                                //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios_ii_processor_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios_ii_processor_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios_ii_processor_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios_ii_processor_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios_ii_processor_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios_ii_processor_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios_ii_processor_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios_ii_processor_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                                 // custom_instruction_master.readra
	);

	proyecto3_system_on_chip_memory on_chip_memory (
		.clk        (clk_clk),                                        //   clk1.clk
		.address    (mm_interconnect_0_on_chip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_on_chip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_on_chip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_on_chip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_on_chip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_on_chip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_on_chip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                 // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)              //       .reset_req
	);

	proyecto3_system_spi spi (
		.clk           (clk_clk),                                           //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                   //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver1_irq),                          //              irq.irq
		.MISO          (spi_io_MISO),                                       //         external.export
		.MOSI          (spi_io_MOSI),                                       //                 .export
		.SCLK          (spi_io_SCLK),                                       //                 .export
		.SS_n          (spi_io_SS_n)                                        //                 .export
	);

	proyecto3_system_timer timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)               //   irq.irq
	);

	proyecto3_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_source_clk_clk                                  (clk_clk),                                                         //                                clk_source_clk.clk
		.nios_ii_processor_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                  // nios_ii_processor_reset_reset_bridge_in_reset.reset
		.nios_ii_processor_data_master_address               (nios_ii_processor_data_master_address),                           //                 nios_ii_processor_data_master.address
		.nios_ii_processor_data_master_waitrequest           (nios_ii_processor_data_master_waitrequest),                       //                                              .waitrequest
		.nios_ii_processor_data_master_byteenable            (nios_ii_processor_data_master_byteenable),                        //                                              .byteenable
		.nios_ii_processor_data_master_read                  (nios_ii_processor_data_master_read),                              //                                              .read
		.nios_ii_processor_data_master_readdata              (nios_ii_processor_data_master_readdata),                          //                                              .readdata
		.nios_ii_processor_data_master_write                 (nios_ii_processor_data_master_write),                             //                                              .write
		.nios_ii_processor_data_master_writedata             (nios_ii_processor_data_master_writedata),                         //                                              .writedata
		.nios_ii_processor_data_master_debugaccess           (nios_ii_processor_data_master_debugaccess),                       //                                              .debugaccess
		.nios_ii_processor_instruction_master_address        (nios_ii_processor_instruction_master_address),                    //          nios_ii_processor_instruction_master.address
		.nios_ii_processor_instruction_master_waitrequest    (nios_ii_processor_instruction_master_waitrequest),                //                                              .waitrequest
		.nios_ii_processor_instruction_master_read           (nios_ii_processor_instruction_master_read),                       //                                              .read
		.nios_ii_processor_instruction_master_readdata       (nios_ii_processor_instruction_master_readdata),                   //                                              .readdata
		.jtag_uart_avalon_jtag_slave_address                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),           //                   jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),             //                                              .write
		.jtag_uart_avalon_jtag_slave_read                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),              //                                              .read
		.jtag_uart_avalon_jtag_slave_readdata                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),          //                                              .readdata
		.jtag_uart_avalon_jtag_slave_writedata               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),         //                                              .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),       //                                              .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),        //                                              .chipselect
		.nios_ii_processor_debug_mem_slave_address           (mm_interconnect_0_nios_ii_processor_debug_mem_slave_address),     //             nios_ii_processor_debug_mem_slave.address
		.nios_ii_processor_debug_mem_slave_write             (mm_interconnect_0_nios_ii_processor_debug_mem_slave_write),       //                                              .write
		.nios_ii_processor_debug_mem_slave_read              (mm_interconnect_0_nios_ii_processor_debug_mem_slave_read),        //                                              .read
		.nios_ii_processor_debug_mem_slave_readdata          (mm_interconnect_0_nios_ii_processor_debug_mem_slave_readdata),    //                                              .readdata
		.nios_ii_processor_debug_mem_slave_writedata         (mm_interconnect_0_nios_ii_processor_debug_mem_slave_writedata),   //                                              .writedata
		.nios_ii_processor_debug_mem_slave_byteenable        (mm_interconnect_0_nios_ii_processor_debug_mem_slave_byteenable),  //                                              .byteenable
		.nios_ii_processor_debug_mem_slave_waitrequest       (mm_interconnect_0_nios_ii_processor_debug_mem_slave_waitrequest), //                                              .waitrequest
		.nios_ii_processor_debug_mem_slave_debugaccess       (mm_interconnect_0_nios_ii_processor_debug_mem_slave_debugaccess), //                                              .debugaccess
		.on_chip_memory_s1_address                           (mm_interconnect_0_on_chip_memory_s1_address),                     //                             on_chip_memory_s1.address
		.on_chip_memory_s1_write                             (mm_interconnect_0_on_chip_memory_s1_write),                       //                                              .write
		.on_chip_memory_s1_readdata                          (mm_interconnect_0_on_chip_memory_s1_readdata),                    //                                              .readdata
		.on_chip_memory_s1_writedata                         (mm_interconnect_0_on_chip_memory_s1_writedata),                   //                                              .writedata
		.on_chip_memory_s1_byteenable                        (mm_interconnect_0_on_chip_memory_s1_byteenable),                  //                                              .byteenable
		.on_chip_memory_s1_chipselect                        (mm_interconnect_0_on_chip_memory_s1_chipselect),                  //                                              .chipselect
		.on_chip_memory_s1_clken                             (mm_interconnect_0_on_chip_memory_s1_clken),                       //                                              .clken
		.spi_spi_control_port_address                        (mm_interconnect_0_spi_spi_control_port_address),                  //                          spi_spi_control_port.address
		.spi_spi_control_port_write                          (mm_interconnect_0_spi_spi_control_port_write),                    //                                              .write
		.spi_spi_control_port_read                           (mm_interconnect_0_spi_spi_control_port_read),                     //                                              .read
		.spi_spi_control_port_readdata                       (mm_interconnect_0_spi_spi_control_port_readdata),                 //                                              .readdata
		.spi_spi_control_port_writedata                      (mm_interconnect_0_spi_spi_control_port_writedata),                //                                              .writedata
		.spi_spi_control_port_chipselect                     (mm_interconnect_0_spi_spi_control_port_chipselect),               //                                              .chipselect
		.timer_s1_address                                    (mm_interconnect_0_timer_s1_address),                              //                                      timer_s1.address
		.timer_s1_write                                      (mm_interconnect_0_timer_s1_write),                                //                                              .write
		.timer_s1_readdata                                   (mm_interconnect_0_timer_s1_readdata),                             //                                              .readdata
		.timer_s1_writedata                                  (mm_interconnect_0_timer_s1_writedata),                            //                                              .writedata
		.timer_s1_chipselect                                 (mm_interconnect_0_timer_s1_chipselect)                            //                                              .chipselect
	);

	proyecto3_system_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (nios_ii_processor_irq_irq)       //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
