��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR���[{�T���CK��TC,���:�
&��d!��]9�'D`�"9 S%�aQ�`!�6������V�W�l�a锦E(�\gC�slu�4U5=1�N�m��l�9ў��P���B�@+yg��=�}|֦���ָJdq�厮2�U�-e�σ�N�_a=ۉ��4L:��^��乥�f]���wߠ/�F{�?��y:� R����E��,=|���HJ$�mR���6v>Z1�o��c01�����'�J�uv'�"q�zL�ˌQbY�6�����w�֮��B�J�� ܟ?��'����
A��O�{z�v�_�Wp3xk,�=����;�Z��M�#c���� ��-5�95D)P4^^I�=��<^?a1-Z��wL��TV��2�n?3g욥����d����K�MX�\.�n����� q:�K$K ��`�#];u �hS�8��?��nD�5M��>3�)��5��2A�dgd��n�~���~W�]s0x]=��V~��;e���օ��ѫX�N϶\b������M��Z���6��l��[��ճ��%��	�ހE����2��ZwI�B���:����� �7m��cJ�J�*�z����9��5�0��)�ŜI/��h9d��g{,ѭ�M�N��*�BaK�+~����5�qʏ~�q��n-��mu��k�W[���r��5�2��^mz�2���x6T�3���M�a�fw0DW�b���uu�ר@	�wS���jy�Z*�x�G�:VB+�2��73��r?��ïp���K��:��<VJ�ʽ.ܳ]r��6U�2��~����Ϯ�5��q[aγ/jy�����m��$�ʖ3������v��5��t�����׋��>F.��� ?���<pHKiP�^���i�l~̝(Z�9E��b�����b���J����D�p�Q-έF������h���2���Ll�-����%��+y�����Oqh����b@��:#�[�J���ÞUə�?%L�P��գ$T�!E�ϭ��WD꣱��	-_ܘ���a��� LeTU��.5o�D}ۇ/#�r0,�0��Xej�5�{�hr�)R�*�0�$�=��-��5�X���z<��D���	A\��+p�\E(�+`�/a�ᰧ��z\�Ӯ�GG����PB������4&�-����U���
�}t�`�X�9u�2j���dk����L��q���dN��|���p-.��K��&��07]��/^���TF!�a>s�C/�<4�ƞo	3�'g!Y��O���B2��ѳF�J�x���Lf»�q�8n��ѥ�~A$~���8q(O1H@Kic_�&J�k*�)��_ -�
Vqµ]�l�n
����y�"Z������M���j�U`b%	c�F�@j�!�h:K_�ʆT�.p�3�`���^Z�;�DS��X�.��2�������W���碳=l	��Go>��vF{N@i��3����3Y1w�ݍ�|�]uO��[�Kvا���]in�`vk�|�Ż�7����$�αs��q��8av��MQ�\�g>W�f���ӿ�:cη���J�%� +�����˲��m�i���ឳ�q6 �aH�B��[�Q˓z0��&t'�%D��3
��o!���C9L9�^�5�c��]Z4<����e^9/�����RP�\v�`���R�ӑi��_D�%�p��[�j�-y����m�����YZFd 0�]��4ێP�;�f2)B5�	o^|M�+�S�=��R�F\EE},�^��L��Y�z
lA�{�����e3M�Ǐ��
j�s�4i֒[��+�Ƀ	x�F�2B��s�NK
(mD�Dn��G ���u'�B:���kw��l-�'S�@ϥ��O�ҷ�ڣU������)�N?7�1���1K�xw �!��_�*�9
�p7\k�i��}2�/3ÁE<�����Eu@���aZW�]��_����#zY�$�R{Ĝ��Bc^Qӗ��	<%�;�z�-�Q�z/��Cc8c���8$����=@��6��ª���V�o��B:�e/��B��vpl�愂���M�[::��+��Ϸ%O��ܳ�th�ⵇu��Ur5��1�Ƈ��_ȿPP��1|C��Zb��~V�ɇ�?\-���'�e�l�#��"9oX}ݣ[�����@�{9�����T��7$AVP40��Z(��T��\T .=�ɣ��|�M�F+�,h������Q���?��~��>z���'yn�H���Jt�h��r�/�}\8�~?0�׻`k��O��hrW4�����JF!m�ޒ� ����m��FսY�H���7qua����V,�����g��2	Kcf�zWG������������m��Z��&���+�_�A�RZqIp2X�B�>d\M�g7:Ҽ�cEe�!���ʘ��>7��f�|�P��=?�}M;0-y߀�}�S��nm"o�ӕ�	��<�$��d�<q�}fc���Lc��vC�K�sw������x��z�%*�R)�]%M�)5�p���M��ΞKn��1S����E���"�>�m��vc�m�F�h�dXC|P[Gk�S;	^L9��=��ܷ1��_In��t�?R�q38K��x�w�HN0�]�jb.��B��n��3�ٖ�i���f��s��g��q�0�V�;�z�(,c�鬘Y*9�b�0�k�Q�o�o��~��AO�K���es�"��o.��uWBA��G-��SΡI#��	BĠ�^ͳq��M!2#�`�P�s6l�b���d���p�IA����=��A�ƚ����DP���S#&�v����R�.)������3o��i���I]���f؀҂I\Q�d�Q/Km����2���-��g��G��K���]�% ]gI{���|eZRS0�C���{�iZ3
ar�_^а��4}�!��z��s��9�@�{���8�ʿ)�����H�3���7�cEva
��x��k��dG�db8<Jj-���]�}m�#���8���@��&1m�S2xy�kڕ[�K^f���p{i �ov���J�������E%P �i�u7��;m(_pϘ�Z��쐳9�,G�?�p����&ԯ����iP������gE�U#�ڪ����hPe�+#������ů�I�N�ђ�ؕ�+���6ꀔ��#�:�����*��f����;t���IoHn���5e�Q�lTq���^/�_>b��������B�a�yF�}����9��eS0v���x�W������'�QQr[B0i�dH�^񼤶!L��#� �So�@Rj<�����>|��/�2�SW3�'���~]�s�j?�x�x�������/�������ͷX1�N�υK�;(�U��/�̍'C����t��;����챠y�꣦t��wR�qq�/�I1яa�!V����q�����7c;A��:53�A^��f��rj%�n
������m�&3��"%=�j���J-퍷�=m�oY�6��6�F�84n*��κ=�h!�s��$��Ils��,�!�2x7k��(���^�&��W_O���R����ɜ3���!h�T�\4��:�Շ�]�8r̤�����VM�jʵ�~-:����P�s��E���j��3;�����av
�"�S��rh5�	b��pxW�{�҃�<f������v�yu�4t��)4xQ�Q���d�};J߭���˿	5���G�kLl�8^�c���~-�(>�G�A�N��28�������;vwCQ��i4 ��)�#��wϜ����š���s�:|�����x� A���>~���zF/o[�x���~�[�q1�9L,˞�wj�>�]ȝ��{$��l;c�1[�!n��@�}
0�|*�ؖ]���vSǢ&XY>�>ㅠ�~�~3��c,2�!��U]=�[�݄��a����+H� Q�$[�c������du�Sݷ�}Q��s\'�U\n�O�ɮ�	��#6����u��p�^/�,�:������k�3'�\!c�fK�H�Q�`��!ںѧ��m�m�Yl��K3���b���]�

!3=�g?����0���i����ك�B�Gm,�*�;"�E�2���N4]�ttA@�9F*�J��!c��X�-���x�ȋh��[۾j0p��ݦr��q� �����ԓ���pN��f��'�ŗ]k��[c!~����ar��"��������m�'<���UD����/���ږ(~u8(q�`nɿ��NˋЮ�����n�X)�����3'»u�Ux�%�l�Sf
������+7��$}���h�n��+R$F_���\<z�ӡ�f����4b���fۂ	�F"�j�s�H�O-y���PW;%B<�}�R�d���Bd?��=@�������׾Ӟ�|(7���ƲfU���e+�1�]E��2����4��f!�����ݝ�R���)��%��*�0�I�qR�����4�eּY�??�<҃�\2B�{��E�sYCL�j�Z���L�kb~�u+ߧ~���o�K��=0�k�ɛ�1�ɤʋnF3�9
�K��[�c��A�;���5=�����k?��|�v�!S���Զ�3����S��2��o�`I$҃�g�#>PQ��~�XkY���L���l�#��`�� ({��.��$7�_��"kc	�,��+�(dqZ&��1Rф�h��I��M׸^�rF�s��ʟ��y��u�����+�q)�{�:�#���@�7*Wu�H	�m]��"92�u�)������B��9D�d`K�'��p���<�O:S._� �4�.�b��0�1=�l��ֺ�����L���3�tN?�a/tȾؚ*efD�@"�@+�^�A\\3��;�V��,O���G\���Y��׌?�	h|!��xz�Uג��H����ٱ]�?��k�A��E!�J��B������ր\3�Ɩ�,���a�K��4��D�M�'{D��j-M���������+Gw+��'��=��]}�䵨�u��{+�2����.���'Y���-M��!�	���w�W��D9�B�] 0)����3ȏ!B���6�����J��AKύLҺ�+���f��>���N�늝BOe���-�l.����Nx+��L;�g\l��L�?l�M�]�䁦�W}