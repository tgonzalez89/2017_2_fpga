��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,�H��#.z����?Ď[>.����Fa�\z����5.}F�?��K^]��WC[ӌV�]��e#n�觔�[����-YQ��rL޿jŨ.� �f�$�W��1�,��B�ֆsv�/nꋽ Jҭs�������7����f���7g��_�aB��5_�Pu�a$ܶf�B(ix�?���&,H�o�������a�k���1����QLWQdX+��v��CK�m8�r�^�4W�y��>j/��__�ȡ������[LL�}b�_m��n��)�' �9�GX����'���ʒ�*¼����VdSY���x�R9)�c)�Uk�s�(P���� &�d\p��D
�#����K����ah� Z؍�0=m�d3S���e��1�I�:s��z3����D��q\h � h���}�{�2�����*��!�₇� ¡�eQ8�R�w�������);G�<��w���b����:�sá9��.6�(}�@�ϔo�p�!Ŷ�	
@dV�v�v���i��	P��H�Dĸ�qrW����������<�컾(Eo;�3�4ֱH�@)��&��3�鎅��v�,[��{O.{Ӛ��ڇCw�vm�^����=ܡ'j��y�Z
��,�|$$A���o��� UB�i` �6��Q����譛D�Lf���k�-��~�l�d7]�����]���]�/�1��?���7�u�~u�9$�M��Z��ш���c��!����5�i��N�=1��=0d�`��ؓ�9n�#=��9l��t�L>ܿ��{S_/5�$WB9��2�ت�գ� it����`��;�����{.�S6��x�6W���f��˚m�~��lY�3�Ks ��v<��4b��![ۼ��L�$�/��7�j�`f���'���v@{�m�E��!�C���Wq\ҷ�0�e�m��r,�Z�A��8R��FUc�c�؍�Q�-FY]Q�BI^�'���.wy�2�v=��2 5�V;�@��Z��rûV��ǹPWyg�1\����sWrV:���~k:���5꫹���z�׆x�F}�2Իn|�9��V�;��Q��`(i�MwǏ���k�����֤tDX���mI��>���է���Wp�#�"�F��똢@�"�2���CWS6-_��h�>be���P	��Ѕޛt�������]��2�����nd$����²a{���=���Ah4�|*2?,�2BA�;}�"�J��|E��)�X�+���'d�t� �}���˒$
��ꇞ�K.qd;��\(�WG�2Kn����
���],h�v���x��ע�h���:���t���PI����s>�ZS���.S���H��-��h>w��+������@���[@5(����~� :��A�iM�W���.}�3|�ߠ�2���I{Ԗ�ӻ.Ϋ�}����ju�]��Ԟ� �T�����6�܄(i��E�\�����ߘ���&.	�x�*�O6���1�+�uG���Z�#JI:�b @~G����b6/>��̲��%֙C�\�-�@����8�Vrg`�G&@@_k68l�Pf��� �s.L]B�ؤ[y�v9.�U/q�E��;�֊�tqo֋����a���!�Ag��3�e��߁㳘����0ژ��x"�"�S$���P�I7��Ɖ�Ǟl��+�"D�Hu�aq��	tݷ0+��B�Mڜ6� �"[��_�� ��B��s�4
L�(�Yp��bδk�֤�]DL�%�-�n4�xD:�� Kl�1��L�X�:ɖNE�ratt̕�×��ìs�R�~���VK�va����Ҹ�N{�9���+k֦�z$n�5}9�:W'�=�|^&:IX�x=3̽d��n�F|U����&옜a��tC%
|S����}���ӌk��Va-��s�N��b��z#I�	���!��f��C�7�כ��!�������0�cp���J�0�Mz�6�aC�d���mH�������~��_#�/��2�7�9�X��ؠ�w%�Ȩ<�7���F�U�as��ML���F,<P��9wT�<��I���0%!��2���G��/6v�g	$�FK�R��9����r8��25�k�`%�m7E�b!K����,��b�v�sk�T�[ĞE�Kt���K�����Шo蝜?h#�4ȼsԊz(��C���N�l��p��ίg�]j�P3/������uO�EqVڼ��I�MϬ��쏄R�Ď�S=�٠�=���ҽ�����O���)�:X��z��j��X��ٲ��Y�!G�Zv��s)�L$D�qJ
H�%�cѾn���P���Jz�M�D�F�Yٮ��DĮ�X��Y�r�6n)s�v-����H�k��t���%��@7E����/�Z�&Qz��ܕձ�uC�79h߃��B�5R>Bv���u�TZ\l�ɜx>�F2��uc�~�:Qۨz��#��Vw2C��w�a�cF��/�<YN��C�eVZ�J){�g(pzƚQ*z�k��7�"� �۵�?�Ŝ���|���"������UT���2��`��BeX�<�z��7D�޼ޚ8fA���S���W�hЁ ���7"B��R�]HS=JV&zIiuR��oE�-� Å�.�e먃j�n	¸�e�!�x���E�q��<�d~cD���l��AWi����mo�eU�O���,�m3f������,�
$�/H��	��jZ��אU�!���FS[a�Ԁ������������5��>��h����7�4MD����`�T�G�"7!�⛻���[��`�d�x �0�`�p�r]�Y�*�����K����b"�N��숳 ܛ�hD���F��@>_<�ne����V�}a��K�®郏[WH�ip�٪��W��r�;�Z��p ��ǹX�N�q������_嚁~�ƅ�H�l�k.E��}�H����@��Pk����K��w�rݣ��!��ċ���t��OU�+��,K��2���8
1�l#m})j�R�� �b,Aly��6�iz�HH̪�In�� �U�I#���Y�&�e�RE�T��)��gv���f�䝐��ήؓ�UT7�z,bl�"eAm�-bZ�Á��?�i�x���������g��h�)x�o4�.������麗#�؋��^�Y�ƞ��}���6�m��$"c8Tim@�(���cm���,h�5�ӶJ˓���C���.�m��_-��a�+j�GP�v��*�蜡e������|\�w��6���;��P�����W�;q��+u[��6ǻ�Y��,�-�l���5$�k�Y5��\Κ4��.�^�(6z06xk@�����J�������H��0��)3�d+O4?���#R &�8z6�G<�����ѝ6T�"\�Q�ҭ�οS��&�5N����,��?5�Xr�RZ��9UQb�X#��&~�B�`�=e(᮸���ơ1-j-�1O�!�����*�Z���*,�)�:��pZ4�x�"��n���_�i�q�V�TV	�lk�V2�x��_��6��!��;�KC�Ca����;\E������ϥ�JPmiw*��^�9Z�L2���yA?�kV��LA[���#��D��]�P�ƀ!EV1$%�dg54��D�W\J7�6N	iܝ+�Zp�Ev��&�b�t��1��!WHBӳ��ؔ�)�wK#��^O�s"�j���$�AYbe��OH&�*e��:A�w0}�}шd�vH�2�C3�T�:D=4��W�|	��h��ޯ�	N����z�攆U�:�S��$*e$�r�ta��.�&_[�}�A�)7��9M��}�+�p���s�r[�#�Qs�R�9��ŀ��~�䴫Ph�I44�ۚpe�������,f�;W���#G7�w��$+,8�B���f�62p�ǭ�	e��{��ADXV���^���+cĂz�sޒ�ޮ E*�2�^�W[+Xǁ�ݐj�cs���I5(dγ�.R�w�Z��/�v��_Z�ɬM"�x���U�0V��L	p�N�7E�D�#RX,߹0ѧW(���1ڇ�$��C�0�;��
���h�3�
��'���fB��:u���� ˆ�PIV���!�o��F(���~���.�=���v��3��ڸgB��)���!GyN�eS���.ϧ��0ج� G�*�Ϩ��yx}-d��/E��fZs6�n�eժ���P�����#���q��Ϲ��s��M���:<��^����������� �����e��G��i�D8j:�"����Z��X��MN�#E�CT�Iy-*]lI�o�����q��cM���EOy��3Vv�׾�ւ��F$��΄��｛������_<�A��J�u�:B�'�gM����mz�|�:�&T��Jj4�`���]z5���avi01t�k^W�Gtl����!�Sr�����#F�������H�l����P��!E���ڴZ���7��ւ��m�:@g��Y��M�02:=l'>��
u�I�� S��e�;o�"��;+�9q:HB�=���N�_M���������(����E��ՏxpR�0�8{�e<]~9-+��Y� (�yӞ�0�X��x��r�����d�?�l3�����I=�K�<���MÌ����d�VkF���s�`������b�o�i�i'B���Q/.{���%�� �dށ����2�HQ��:P�?8͒������5)�e�l���Z;�����qfjSW���:��Jw��\�oֆX��#���x�+׏�5,��Z����y�ϝ^:��1��EN��ݤz�`���r��Y00X�s��6�������}������#�C:�hk�"�]|毎°Q��V.R�1�(��q����&e��;m����:�,���Ny�G�sNe�\|�@�C9�閖9��*�[̅����TN8&���x	��ŭ�2#��$��Ak���%G3H�A
h�r�LK2���G5�1C<1sl�	�Y?�935���ኖ�NAu�Nv���>��{����N���K6�A�.B{*�x˲&�5J~�fɭ��"��� �8i�"0�F,�u ��#b��`��۵�S���
�mW��|$"��q��]�咀wjj�i[k����}=`�2�	V���^��3"�������l��6�Ƕ�ũW�
��ݒ	ȿ*2����/�)tq=Sx����UE���O�[׹��+���>�.%��g1��>���I�Ɛ�S�QM�x`hV�
���3h��9��%���y��S��p�j��H�C���W���^�,fhK�� �T6@�����]c�	1�-���6���\�W#�ni�̗���[�BI��b��[+��X<rJ�4�xi��jX�>j���ME:g�SI����QK�p�:7M׎�_&,��U�!D��s��cW��d�O�-��B�m�(�k�� 
�ɚڭ�4�����U��r���08�4b��h�f�wě���c� -Ģ��H�������I!}�8�(�5��V�h�qW!;��̈�����Ǣ��M�� lR��D%���<զ�ޅ*�KG��CϾ�T0�2]�Qdϵh��?O7��X��\��[�n���힨cS��1�9B�z�=�)�~�	�^�Bf���!�2����!��s��<��k����HG�����Nx����zY��-O��;����w-�v�ּ�F�:A˅�8������ի�t��S�/�s�6%��|`���u˅���x�~��xX�>!��9iD��8�o���B ���u�;cs}�C��1���r�a�x����*F)+��%���1_��3�*�8���m����p�W?�����._��P޺^*~��l�<��V �(�7aɽ�e�@�n5{��t�X�Si�ȅ.��+<$�჊��8�c��Y�@0I�yz���f�ppȞJ1��X@4�̜�X<��Be 6�
w� ���l�v:f�%��N}������:^�.�o�M2�\B���������aR�@�;�q�2��ݨ=���)V�AP���&��$>깥HS���⯩"�'bbK�ah�_�g�+qE	ʱW3��l+|B�_NNͮ� I�e�{sSJNӊ��
�����G8��#5�k�f8�.�!��>rPJ	'i%�����%?E�Ln/�Lv;���s�;^�W�J�s{}��89M?XKZx>=r9"ܫ,�2zy���-ڍ������-����
�s*&����}�IQ���ףʕ<�o���g���J��U���Ւ����Ѳn�x��#�p�UKF<����h��D� �0�;42�|��
�R"Gtk�&6�vƷ�Lk�իsb�M0s�����菹�D.����� ��BJ�X�ɤ��a_��^����`��D���i(/��
��a�$�s�R�zS$s/Z�L�~D�]����Fl�ۛ��S)�ߏ�K�A�%[d� �l �dH����j"���y�r��+h������P���](xͽp��W�v�V��JSԑźxYN�Z����f��!F�nk�V���xT�R=���ni�w����O`�*%EsM�����S�,���"���A�2:�*��F�4�]s@�%�M����>:w3�	+��?d�rH'��jIxq"���g:����G�64C�/ݸ��Mv�RJ�753��%�;$�I�S�k�����k�����IQ>4wn�en;�����D.����p��<�)t�Nj�,�%�lwLM6��RE��{�t���(/# �EyH*
��FlM��c{�u%��I�8d�خF��S�136���������)L��Hg/��F����4�3U�B폊{J�e
�� fJY��>?�ٱ���B�V�4��u���t)��1�������l����˖�>�ƴ��uQ���� �o�^�Ic0�;��ʜAV���1���<������0��a�X�"7�������'������$�V�o��Y�3�z��Ȉ���(�:"�gE�`#�j.!%0� )p.���z:�"�	�:���Ɵ���O.����K���6�%�uܡ�Z?�E�I
۟c>
O¥qg��b&y�f�C;rr�bJI�B$�i����M����I�#o�)�~��"���f�������Iw�$�>��Y	9ݪ�1�z2�O�x����G�fd� ���˔���lu4'�7ʥ¿����DI5:*�db��z`���g�M�?��r����C�^�B�70�F4�|�s���H�`�	J,��z�T��S3 +��15�o�(j���~G8�c�cg�!@/�	��Ω��*K�q���J�|��O�[��Au�w��Ųj+��伔���H�)C&��~���ښ�}�f?�Q
���ʑ��;.~R�S����UD����tQm�����d]�����Rd1���S�U!����сZ�r[��N] ŷ͓��+T���Sj@��!:�ϕ��@��	�pqc�{���U!�e����{��wi�:�TH�B/�xfxv�_#���� ,���ƫ���y`7x�Mm6�s<&�`}2�d!��=b!��>�
a���w9��� "�N�3T^���:Plw%���G���Y���(���6i�a�Y>����$pӎ�u�Med��0`Qh��^~�o���o�3����ڢ�ֲX�ȟH;�M!!�`
�\x�/��Vbe�-����bf��z��\�8B��ӑO�%m'gm���l#��X�%CbQb��@���pIZ��K�B���|��7�L�'��&�@���Q	V��.��G�Q]P��4{��B�9c�f7���������#��������?�9�Fw�?�PI\^�*�N���)�E�}&��pS��N鐨���Qߞ�h�s]�2�{��lV���
�Y�E�F�Z�u���eg��[xbX��b��MW���5�ZXɬ����w`r��讠OY>��2�sM�n-�S��Z,y}��� ��pȝ��.wb .)�I��Dd@{G�Wh��	�lŠ �n*�����~r�NvBu׬�C���Z�pU�*�y�9/|��[(&�Օ{
�@lF_,/x3m*�"��p�ed����M����(��)��A��޶Z�D9�� |`$O~�� �!�>W�4뾈XZ�S�]�	.lT�6��L�"�]#p./
����f<�:K7��$�+�����xC�=,I������=�u7<��z"p��\xy�8^�nL�ɮ�B!� V=�37���{0�RBd�?}����n?;B�1�������xFL�ǃ����'ܣ�\�)g���9�14H��;7���?:j��E�ltL��Q_���i���uq�D���>UtTTT�t�܀:=���LÑ��-�NɊ�/آA�Q��0��I#`K ݉6����%� Ț_�b;6����F\��R�|�+Rr�y��C���4i,R�e���՗̉����5���:\i��L�,�C���ꈉb㣪Y��e�r�Bػ�wUE-���z.�0��8� ��|B�ԁKz��N��2#���HG:��6�.�,��mH:��	un��!��5�D���H���$���}�f������(:�!v\?��dP(k��l�=Urx��^q�$�Z�Q�+��П�]ye��!^�%T�Us"��d�p9NQ�|��H��Ld�%Z�N�Lh���3�Q������Q��c�T�e���%�R�\��F�U(:j��E��(GO� t��+6��n3��2>6r�;����%�%}C1��>�a��x��� ��"�ȱ&��$�]��ʛ����	n�j�Pθ�V���-�
i�ī|bh��}l�'�zkQj�!}gG�g�d!�RktV�����蓓*A^��I�7���\�o�o�g�����X٨q��e�z�E.g����(�L� R�ۼ��F���o_��d.Z�h���
�OF�9Xz�(2�H���	M���K4����X-�l �y�%�(vF�
��Z�0�D^�ph��������<�r�#V���?���&���� uN �ҍNZ�S;�MS�g�|.}��P��J+c��Ub𺄻�6��B����t��s��ԉl����a R��kT�%|�%`nr�����i��;�ڌ��y�p���rӌ�W4"�\���@��M�Џ�Y��A���*����f�&�R���KtW�
��Y�]�W����0m��@H=�${e,ٻ|x����[�=ٕO �>/���&�4�w�V=f��E�+.����˕�-�A[n9_�u8�jxJ�m����9D�b�2�%�C�������Z\�t��]O�4�G�_�t���fهD��U%0l�D�ƐɍEX��:�.�B���e�3�O��̿;NE�8F&�?&��5���_moM��a��l��R��> cM�md:H�x��q�|�>8�>�J�t��f�Z�N�[̏k,e֏����p���(K�7F�&U�
Ï����i4ڧ|B�q�@R}}�e7��e"\_�݁�a��l��N
�xs^��A.ܡ���3��%�[g���oSa��>+���b�S�)���"��~��%���=��� Rq�pXw���!������q�0q����e��ؓ��U ����m����q��\FMMfzY��3���d���ʎ�¾m�A�-�c��}[�b�d��a�r- T�a�C��!c �����@.Rğ�L�P��I�x�S~���:���s��e�"XI�l�>bw���u#8���[2���(0V�i�޶��H虌��%E!0�_:��"٦s~Y7�h����?&�v��<��'"��=9zۣ� p�R���)뙓`��-oȐ�iF$T���&��?ٌ'�=���I�N���P��D��� i����� y�(?L��Y�t`Á����π5B�.ß�)��\����
�����!��E>�m�Z�	UP�6��/�k��	P��\aC��`�A)+��Űls����$�-�-aj����&�j�R� Dht��[�����$� ��SD�ȧ�=��J��;�e��3@!�I6�0Ք�t��F���2/�䓝���l�%9&�-ް�++U1���>��n����#Z���\J09���Ꞩ�uu�D�(���be芣B�;j��e�3�F��z�?����;��ū.a5��0��UX
e�s7�'r��j���O��!FPE�G�Xf����Av��]68o�O��96� V=V�n��	3>s>|y�3b'K)x�5W�o�D�Z���!�x��٬�%���������ζg�n��JH)�D�o�}�l)���!x{4��i�㪅.��`P��i�L�)�8��.��һԒy~դ��O}����@3�^�$8�c^,��A��e]1�q>r�"e�]�di �1�Ҩؽ�z���J�>s���-�U$��i�>m貗}�-�^���+����`A�
*Z���0J�q]�. �A���w�0´z?�?�^%x���Mz@���l t e|Gۉ[F�7ry(�4p�6�H�B;�bYZ���oYx���Ցg�;�4p]��D1��:��٫?�3�a��se��0���3�ZK��є�5t�>U�q�Y����� i=v+�9+�VKq̺k��L�?��I$a���*
Ieܞ� v@��6p�˃"����_qz���2?�Ӯ���$ۿ\|�R.�C����K����������lq V���%���b�L��u����]ێq�o�y�j)�I��L"s.ݾ�&3�y�l����J��T�|n"�
�B#��a�N |G�I��� s�0c������oO���j�ɩ)�.j�ލuP^�v�x������굆��Iљ.��D�9�����}h���(�>Io��2���PH�v�N�1��ET*Cb�$8��ڽ]k� �N�%�͢�9�7�Q� e��v��Iu%i6��G�0�y�f�{���(�o9�ͥEr���J85cN�ưwA���1����VL���S׊!�u_��9@�)H�B|�T��?�j�e�ߺ��@�&x\��v�TWׄ���%�8U򵻩V0�ێ�z�֘��*�Ą�E�����mD#�$[jo�':�Nl4G�O&�zV�t���ܫ�i� 狢}�%��Z.����{��r�rtl&�V��L��U�V�?߁��Y�9M���E[͕rU�2f�7?d�=��є�ղ����EѪɱإ��d~Z �����$,9��S����r`�O�4�_��{+_��5B��[@�5��2Lۼ�����@��n't�m�1�sB��W?~��F�-O����]�<]/n��	*B&PP+=]�=L���WƐ��1X4m�U������ ×m��K�F͸�����X�$�]j�v�z�F�XD�k:�~��YIIe!-�d��b�س����B>��%^�:S���0����ȥ%��XY�M�w�\}�5�|�s}�+�j$[�$��n8Da��9´�{�l3$�E��9�ŀa���<2�PPǨ�����ݦ�!�O$��j9)�*՗]��xJF8@�2J�(����v%j��Y��`�a�x��
斊n���HO��>�*`=ubbdbwz��i!TP�<�iF-��U�����'����Ou��f��f<O��������K�E����l'�;v��,wɮ�yvᕨS{�����nO��h����o�U�H�R���geS��c��u����tL���5-����`l�3i�r�΄=n�[��AW����	�^�΂�U�_�{i�&�_��z7I/�?b�K��RAH7n��8C���S�%��ة.s6�'҈g+��V� ���T�|IdTw����54�6AT?m��ڤJ�&��:�k!�Xf�룧Zp��k��{��+��A��)�� �ӓ2�T��%e;����=8��Y�'K9��T��f��fWg2w�tso��D�yik���<��b�)_Ϸ,���dGq:��Ϝ"D@����To(��j�B5<���$T�w�����S)��Rx�Uկ
��Ӭ&:<Y(21��2
_@W�!�9؝��/�vgbxxii��՚Or��
(�Zǡr$FX[�}��/r�ڕg�z뉄۲=2#L%��Uc����0Do�"�?4�|�(�Z����c���S�*a��=v���|9k�
/ ���iz���Vn k3A{r��:bm�x��E����T�8yvd�#�AN����]��"�9���d^�T�,qq���d�c��/W"OH�������!��f�F�1B�>	n�¿�&	#��]P�=�K��������5��S���JI�r֡������ov��r"}đ���#З��ر٣�̊��-��D�D"6��C�S�k��h�p��	������MVٺFGȰ����
'�ݜ��ɀ)9�J��AK:?ם Q� $�����D���V���&�܍�OK۪��x�jΧ��{};�=5�8m�����е~I���rwIA���
�ag �"E��Q/�H�p�����lr=��3��:���w	>���崙���i���Px'����3<�P�2�-_�r�H5�dL�-��0jW�XW^��i�xQ�@�F���6Ce6U�缥�"��k��<ˠ��&���\{�ڵ?���Ҁ�G�N�BFk�瘬]G�~r��@����d�Jw4�/�VS�4\ВPl3 ����AP>m̀OQO%��U㨒�\�)���� ��%�mlB;o�閾"i&^�P2��*��]���5xB_{�k@��22����!��W���9�.7���ĵ�t��KD�F*���2��a�z�kKݽ�DMyD�%�}D�)A�'ё��I�>Γ*��xISa�CC�'�TB��	~a�c�?�񡃆�,B�^��G��jmL�
x[��"��߁ �f �����=&c�����������!�����Y��f,�{��b"d9����2���R�%%fc �5��� ,`)pԯ���,7{���I�*	3�m=3tk����ْ� �~g�1pwk��/�l�j��'����W���(ɐ0W�m� 	,xe�����Yhդ_�IK��&���^V#��4=Ss2����Rv�X������f kCY˥������}~�=w(�!s�?����p��7s�d�p��^ �q�X/#�jʑ��ޝ��nł�7 r�(#���
�H� N�'$t	t>a/�iP����Ѽ����J���ap��ɪ#�߂;�g��Q��m�6?�݋%��7���h�3ޘ�O&���q[�(+�wB}'˚�+kC�W[Ѱ�)�J�D��1<E�1w}��C.?B� X�i���Ek3��w�Y7PIN�[�T�N+^Y���X����#h+�1pZ�6�i]�Y�	���=6tD�B�S�����5��9'�IJ4w[���5#]=�&�n�6���q~���<u�aG�C�Va�ύ�	%�_\�ԙ��i0w��|�EgU� ��-�~U����;Xؖ�%������3�� ���ӣD)e�؀A�9-.<5����4K+3��eci����@�dw�o�����c����b�A��jjΠ�L�C�3��a��t�*7"�~�!|�����=���V&���#F��?^�͢��O��'sC�H^D�H�^$�]�n�sOj�r��Q��#�O;��� I����]�f�6��X�#�fƼ������I=��k�����V'���Ő�-3�jy*P���������oO㷙��Gr�7��pEcL���>��!�9H���c�uS�L৶k/HT]��Z�~6�=���W���Ӿ����.��S�:���M&2`!�d^���M�v��Z�u:'����x>��ۿ+��U(9�W������D|ᐖ2�(��h��� ��`��}�h�9����~c���f�U�ư�h�C~���О�Dk��j�̍7��,���jO��ۉ����Cܬ�ctL�O{����h/�o2/QUo��u!�4M����^h�j$t�𪤖U�NO^ZH�ѿYf4͘��W{־����]�ʨ�6z����w�`z�e����+"��c�Af�g^@�hy��њ�Y��r +���}��^�"aE��*Hh[�
�G�
�~?鎨�s���
Uk���bm�@�{���;0�}$��� =��$%���	_"�E��=bȴ|��s���(�:[���.yǳN�7�U�( ��>:
�^��,���r|@�	y�x�~!t�jp���ا�l���ߣ-͏�h��K�]�{)r@=�~O�<����r*07A�e�F�1&؇v����Ԉ�B.�=u�'����\��lJXH��mw�y����	����s���������9.Wv��uN�bR�>�}�,T�<��bDXr1�hCR�u\�#��0�gs ����^��7N�>�*λ��@�_�v�h�U}�����f��H�(:AT�`�'ѥ=��l6��!5�#�9�C���e�5>D%��dڰ��ٷo�����k�
L)�Y���%�[��T4
���ZrO� �+;߿�\�ˉHF�UV���߆��j�����Y�	��6R��ϰ�}K4��g��Q�̯�G�K��WzZ��ӝ>�V�� ?i~O.�D말j#n�i����/mFL�jwo4QJP~�Hi�g��|��5O�z�5��m�B�n*�.���D���	-�J'��8�%�`<�8��2�ut�u�w�.%3B�UzS�J��-r��'����Nq�����鱮��0u��T�};U�	!�C��3�U�#K��RUSȱ�b�a�4a��>'&���q!ĺY&����u�B�-��bfC7-���=�4S!K�$���-n�A��v��F�����kg��zQs����"v��ge���A.c�Z����plt�-*J�N}���Ux	t1;�?��cv�H(B�� ~�/ �0�؂��{�����"�C�5�t�<��	��Tg@e����jv��FW�R7���:�e�]�Qp�Vn �`���8q�����q�8��+A����;���<�*G�Fдo�E^6T2K^}�y�{���}p���O���R�>Yhf�*��-E��� AǍ��z�# Q�s$>ޜ L����Y�7,��$.����7iBbA�����%m�ȸ�[D��:t��z1 ��k>�zhkm�]I1����W�*�zf����9��U�TP+_��-�������t�U�ioߑJ瓜�c����S�s:���?cj5&�}�p�}Ď��7�L����Ru#��G�]D����B��g�&�%t��i�x�c�٫�,�Lrd��� I���%�x/l����Ac�`������!,���z"C�a=+����b���hw�Ӷ�`r��(��	�Ci��w�
�C�oz�������߰��Px�wvpY�ds��>*�{S�X��{
K�V��Wv��1��?����Fhȝ���H���J�V|�3UK8~�&�i�輛���:�#>��4A��	
Y�d��h�H�����@W��N��D��$����e��rU�{����"��dY<�W�!��������=k5�:?E*��\=v=:B�ƍ�D�!k�e�8sݐUfMA@��	�sI�����.��u�ׇ���O����G��ul�z�u,�	.T�"��w�0��L��2O������� �>AIU%���PH�,u<�|b<��Y(t�f���,����߸T�F��<Ȇ,���3��{�:!,��y��*6��աV��i�A����o߻ ��dof�a��g4���L�3�7+��=O�O+��,�u�d��8��2&$
K����^��G��V���P���zx:��^Ɏ_^*�&-�D.j�w���s��Z�C��1dN���3A:T w-�7#��؅4���#0( ��0�FQ?�b��:T*ةVc𔞃a�ӿϠ"f�,o��"�sy�Y�[�G�?�b�j?���^8
�q�����U��PRk�{?�{�H�E�28'�޹��ᾊIɒ?��)w��-�B��r�*�OV���uސp�>o�g���j�xiӸ����N��k�-ib�\�8�h6s�&�]�Ph�h��D�'Yx�|��!�܏�z�2�т?�D֩��xՅ��㵂��.�m�Iץ�@��@�Q��Ֆ{D�t����?�4%����Ȕx����nE���t7�j�X~z׶�Un�0���C��t������rοo$s�ÿ��N������G!a�M�w���,13��%+'��7���R���E���0�QeY��f��<�YH��}����tX��H��)���� ��="��+ɠ��kn�t��r'��%������9LSB��
�c�J3��T%���]*������cvHcYS�$��;�U_��<t+� ���8�/ν]�b��`C�� f���B�������i4��H�qa���u�,9�J�LՐ�Pkux3�E잗b��L�`DzT�U�<�A��FJ�BC=p�X��KNE�T��6�� �a�n;}M�96��D��V����E�{#��ӄ2� ~)c�\5zb^3�(�+gj��������e���iU'L���c�5��+底���c&��D9�w
/	��~���x�4�x�I�0�B�˰h�Vԛ����F}��`�kf���:T��t t�xGq���j���e�h��X���L�e	�ܕ\P@�1�j�7��  ���C��X�������Uf �4:��+s��8�/�~����GVT��5�%"���f��~�������%V΄t.V�5I�vAH��a�X;9&�����{��Wo����8pT���{�]��B90����Eږ����S�\����B�9��O�T�#d�⾎��j��x���^�lwԽ#"���֘u�V��%�����<��"�X"��+3������!�^�ڽG�������[:�}�_@���7ll�������^���_ä�$2ӟ��I6&LO�)]}o��l$�{��ny{�
BIP79dET�2[r;�{��fp��`빘�*gw�<?I��F���#!���<Bn�?4'ء��F���e�,�<xŴ<�`��%���:���j�VR���N- ��@o��iLNF��o�C��Wދ-	f��!�6|���K�Q��t� ?H��S>z��Ä���|��c3��[��3L��h�X�>X����V��+q�:G�d{"��
uh����}aO�2��\�Ws��$�C�7>�:���'��QWd�wmM�|��*�w3�xZ�����Ю�����@U��)9�v�G����q��#��O���QxƑ:m>:�FW]�5K?�CPr�D�dt硩���8=Se��f��2�l�Ei^Q�g�A}s+��T�g��^�A�q{[���,;����~:[5bѼrHm��Y���._�H�o�D��l�-kxÓi0�T+j:o,j��&�QAS6<���f��Y�7�՗��d��
��`�#D&��D�X��C2���A���f���$	�i�L�m��Җ��p�W��§�A�j�nNA��
��˒	
��Q�S��Y�� B[K%�iV_N�� ���m��+��K.@�.�.�2�XtJ�,�-�k���h��=Ȕy���h��e! j�ć����zt�g͞�	�ͫd���֪����_ ����1m?���+F�;�t�7��c�!��T3ڲ�SE7;�͠�!�lv�y%��qq��� <�XEr}�Q8�i�4.U:�j{wXE�ZǴ� b_�3����TR�	[��Y�D��]J�1���j��$E
�6ɜ�Y�a��Bߓ���(����w��h�x�I�77�L4(YR��|�p�=�@ � �5&���(5|�EN��}o�(Rq㼏�k�	nG�"�c�1��GN'X������|�/���G#7tp����_�H�
6:��ys+����<�b��YH\����������ua!,x�W7}����������Jd���Y�~o�CoGT�g�j�"�#5��<��&e��`��G0LT���]2ڣc���B��_f��[
�E� r�'
�q��bS�����&��5�2��� 	�����u]���M��ݧ����)�����t��j��}��C�w^V�K,��$9Rz�����hЀ�O�����Pƒ��<�6�%�FS�bK��!a�䯚��� g��lW���)�N��g��J"Q��2�B��+N^��Xi�����Q(4�\ە7�,�w�oQ���I�ZN22���6��}҇��ѩ�V��#�h#��:� )D�d�;>g����9����\*��|����XbV;Ʋ%�5���GMAF�qJh�X�5I2.+��b
��Y��;,Z�XΤ4�"������S622QM�t�dr�#_�]����ż����|+�||dĪfN$y��Z��]FQ\����tG}BO/*~,͌���7c�;2ۑ������>3�xL��N���eE)���jy�AԘB#C�kף��[=VgEB�[��\*��J&n��59{TR�2���-q�mM��n�S��Z�n.��_��^��Q���O����gvK����'}�݄��pq��haT�G$�/��'��h������u����!R��X%^�-k�+�FǞ{��t_y#�
��D)���Ope׍\�nZ��%���]��!bj�f�9'�k�&/
U�S�k����u#��mL��Wf�ٚ���c�_y/+����,�
_����(�/��\����8�ܗ{��m�z]�-0\;,�˾Tu`�PN@�����i׾���,B<��ih^\�5Y���@�0�:����@�Lj���r/����r��0�ɰ pq�����E��ܝ�o�	^zXҏ����l+cEsb)_�� �b-v̊�J/w����%$�eB��gYm:�$@@I�aA�7(��t�-�
o�Vj��j`S\9(�OV8�{��S�l_�P�=Zibj��[	�49�1�W�_)Z�L�JBph��AzFo	��{���cEf7� ��:�c[�}fh��398;�c\�h�p{����C��������֘W	�۾�OU&κ�l�ʑO�W ��p�\B�
���"�t���''$��% �W��R����n��Y�P�;h��%L���
n�mt�JO�3��9j�	�*��f��8��t+
�CD���=P�z1��p��yp�����h����Cb���b�~~�Պ��G&\7�;ĕ-P���!6RC����"�����K�3Ѯ,A�V-=�R��S��H�X��d[���Ɍ���ݧ�'��}>�h1T�.�Hn�䱻>�0�:<���"L�[8���m�SCx��~L���"tb���T����y?�'PEƼ?Ϋ������mcEБ�����=��?F�>)��|8~�'��<��]
�Ha|/4T)"3a�}�N�da��#���v&��lP\��1Q���W���zI��<�}�Lw�ՠq��G��;����h�Q'��l@�Q�n�
ꁖtΫ�@>�7�-V	�����6*��	(�V���> IR�`C�H37��C�M��`��\��0�6{�9bE� l��e��k�� `f���}c�敉�����#��RD+�\{��1�t�gp��Qn�D��;L�ᤉ�i�_CH�%���|3�懶�aR�($5�O�#w��y��]?Y�(�
ԕQ��f�\@x��v��\�F%Y|e��	�F�,���zN���Q�g�v�u���4��t�5�<����sj���,��Z�bN\���7�O������5�(����5C�)�8�r�i�:y�EU
���:�W$fQ���ae�a�dJ����%-�)����Y���g,�Ύ����79M��Q.�������k;)JA��F&��<���H�ϐܓ́i�84��,����zTՒѭ�o�mʐB$���|�@�:ṧ�n��uj��x6x[���d8�\�3��m�.�-���.�' ��-b���+�A~M���ǫ4�������Rn��gg��cv�u�,����~Pz�^��AAęȑ�U?s�H7~�5�_���un���L�8�Ȼ�)�k���de�^�����ٹ֑i��G����E�S��,�9��z����[���\Ei݄���kjmk��b��i@<�x|�1iԍ��q��K����-����R q��ɇ�J(#AC"ٶ�*�F��C!1ִ��D��6�{f ��oMv�����!��4��P�=��_@�dh�����s�X���H*����>�s����nXReY����2����Jaݠ0V��D RD'�xW.��T
�`Օؚ$�����9���nr�����T��\3ԣ�C���/���97ftI5Dߜ|�-�K@����S�}C�ީ����="��g��ͅ�Ė�Ny���nOC�rɫ� �.t4+�T��ۂ�aA��5$�eL��"XyU���UG4�o�U��??޿t򀖷���|��f�n�2���.�?����7KH��s�M��h�S�S��?��,p�dQ"�ǹ�1T��3T������_�Գ��|W�8-��rʁ/'"��b�d��Yn	-����%��s�hf ��1%l��pa����!V�ƕ�p�f*��h%���ؐƙ"�9���x�vׯO�`�cN�Q�[�؆G�����D!p��|���a�Ok���ߊ����5ƬD�M��9�����&�I��;���&��"¦s�PҠF@��]�Q�v,��;N{}���#"ƬD�ŀ���q���oBQ��<�	���;(y+䪚W7MQ��0��|Z4��V���t n}p��3O1#K��t,����K�F41丩���Kk��t@e�W��}�������n�\Z�5�)[�'vڦ\"�;fP3ȺPH
D�եO$�{gD��z��:�Ԟ���I��溬tR�u�d/=�|�rR5Ź�6��D�C�0N��@�K`|��-�gd�����pp��1ָ���C?ݦ�n<�8��p��j̋G� ��x�zG�;p�d.d�Q�n��^���T+v���Em&c%BObΗ�!�\`��y�$��`��.6���4�=�*f6����ct� �n���0����p�;��"E�Hjfg�ю�G_xY�.aě �_��0A��1�G�ہwM�^��d��|��Sqb��0?S�P�I�1w�
��~�W�
�o=~���^���������;�>=ypO����Ω�㰬��7k�k_a2�5�Z�Ц�
��:�Nw���k���@��^�]k�7�� ,ӑ��Wz�D,�k��ޛ�dXL��e�!�{�O�?��#a)7Rr�%�H����b4:V�9@�G�mM<~�6�7d�:���~�SaC�A�a�� �k�5O��A=�>_���w�����h����I��g`�VA���{�9U^T��tV�9�k�P�뎽w��Ɗ���3i� ���1h�w��i8�S�p�u�Kn��I�v{��{DJ�ťc)���J"͏|.H+qfL�	��ȉo:��>
�h_X^r�!6]!8��}D��HFD�u\����P��+���7np[�J:��S�Ę�=u}��m��N�	[:}�ŕ�Ō��S�S?�	�Ǩ�n��LHZ�J
�u�Z<�6��Z"�R?�������uhsȅ�H��DS�Ĭ=��6�샑O��-�N"���ͫ���Ii������� �F��J�#���Ğ�5炽6:��'�w��&]��H6�%�����%��3�P0�'�#������qNa�@w��)�I"vd��7�%��}֑�2�/�P���?'X���KZu�-zUn=`n�WZ�Ԅ�I�4�[���� �����B��`c������}���X��v�ؼ���=��"��P��d�Q'��=�m@��D�ML՛5�� &�hf��|�;��#��&ߕ�7Vp��{��)狛b�e�;�Z7]�#�7ڏ6�o3)ꗿb�~��X�Ӵ�����5Ӳ��U������]�YM�xi����@����������{;�U���{V�}�=`l
��Җ*�A�{�\D��V���-�>=f�)4�s2z��aM�`�PD|�B�����u�� ���
��4�3�͒˅�*�R/o��Yx�I�T�:܁�=b6�<�*�]�
4(��U����ŀ�f�����A�1ZkS�\�K@gU/=P�җ�w�Wu�{lS8���
rJ����<�Q`�P`W��bL��5i��7���G�6�L�:�6)q0y� �ۯ<���C²����	����jBDH�Sث3O�]���,�\y�.({!���χݬ�cы?�=��4�9�={�b�
��x��%g�N$}���3�TFZ9S���ɨ�SƯ�����~�3?�"^[F3Y�J�63,2�!�E�s�5���[�Y�g�YbLE�'�:>h�	�Z����z�3�n�@�z�	o+������_�]x����x�V�;���LRV!����W�y��ů�Ȱؾ����|R�7|�{v��[������6�
�d���>z\MIO�f�079d�U$�,�x;��(7Z>뫜> ^n�����o������ <����k��=��е(
� �"���ƶ��M?�ɾܓ�	�ĝS7�ꃹ�0��R�-��c�Ɓ���FR�dKT��ӂ؍[�)a��;t�Hg�s\�T��g�����+���T������Q%����W[3j��y�����4�ӎ�]�1����z1�D %OJ�|����_��|��+�tǥ�3h�dPb
S0��3�Y��aa#o'}�J$H�	#%3���kX�!ZB.�i��	�V���+f��H�8ۉ�d�f�db�a���g���tR�Us��y�|�3��0����>�=k���'��WF�FOʂ}��3�--�i�{0>��C����4Ý����d�P��~=GA^I~>�s�����3>�ɏ{�#
K>M���.Ǫ���0�ݜ�Wg�m�F}!����1jLbW�Å���8��.z���]Գ���w��қB����%��.@����JgM^��/��>�Bg;�PJ�g�}lO{���Bn�N��1Ma8�F@����75��4���RQ��*�2:��=
(W�o���Fjɾ��YF�0xUjc� C��������c��Xğj1�F��b�ӛ��S�S��� É���+��+
h2�3J�)ʟn�o����DC�>{_zeHHS'��&,pR����hH��3��R#4���V0��+�QE�`�<��PW*��C}��=��y��Y�
�R�u��e�~o�Y$)�,�
*��Q���To�Cǟ�z�����_%n���3l���w�m�J\W.��Sk���ɾAP2�ܭb	Y�h!�|��&~I�O�X>M�Bi�9�^C��z����3Ċ_lI�~=�Q^`��>v�NtȔ֮��%�B8 z�;�<}J�>g2iTkg%�9�T��`к؜s��\��]�ꗏj-��KSϱ> Fjd�lX�dJ�
	��X�v���#n�Z��ZĽ�d<������EM(�M(�:_Nsת��B�11���;j�;}�3ꂫ=�36�  � ���o5r����C>H��G�q� �F���ri�^���Ç���~�����"���̛^��F([��Q{p�]!
��+h�g��xR!�S�9�zoZ��1'�?3��� ���\ʀk͠�!�`R�|���x���a��0i,.���\�8��i�or�~t�(�[8���AQh2�:0�rq�<h�vu�N�wc��[�TR�)�>,W��jl��?|#S���D�o�c����U7��59ŘQ�t�$>��^�v�B�$kY�R�p1�F��v�v=S6[0��a����}��S�[=�dm �S� ��5jO=C����%fV�ͻA���dem�0:*G1���-���b�
�t�o�K�nM���!��k��cg�ԗώ$���	Gt}|��J��T�������� ���ǿ�m�C�LD��Hf���MG-�<i��������ױI�y�ߣ�σ�HF��I(�����lӥ��f ��^w�{�nċ�l�.< &�`�/�W~I���*��"YG`Z��TAݣ�:�$h��6!4��թ�e�Jl���a��ц��VJ��W-�U�.���1��8X0`'��g���f�)��?1����H+$���z)��m���Ms��-�����F�$����_Ր6ѵ�#�`?:��M�Y��vlY��W���̘�[��,m��B� ���殜omc�/W���#+��f�1�Y�Cw�@f��k�1�6O�ꃉ��J���?�Hg���P��/*=���8���hu��\�"��YI@\��2%'g�\�����桃�)�W�s���)�R�Q�kh�(�W1gD����|�����u�@�U=�۪W/�+�<��T!��g����V24�U"�$��f�.J���%�֨±��Ob��A��,��$r�zv�H�;��^��f?�0�5��;"
<�=�{w,��?�~ Q����@���д��X��/�$�f�e�?��X9�|������u�Ӥ'�g>LJ}��;��� 9��i9�4�1t����n�}&߹(p_"�ͱ��tX�=��<�`T(޽�S�l��#�A�~���w� YV��fKT�M��̇$�����4���[�ŋ�_3g��JV2�u� $��2|��h�Xm��OjR�R�ݯ�6��QA���y�W+��,Rv�靌9�9�Z��}v�N����ٮ@2�/f�"�tyͻ�G -D�)@��+k
�f�+�ݑWO�M�.���:���X��/�[���w�@���<m�K��i&Y��k��|��WE�;h�KJ����sl,5��#s.���2C=���DĽ.x
@�K�SN���]'P~��=?%I5W5�<>��;|!�6"϶������>�4�'Yz}��	v�i��Sn<>�C�Ms��S�
ho��P`e%�ǵ�����G2��D&���qԎ����#dTi����;<����=�Xܱ��XhGDP�Ph�-� ��T���<���d��g_�-Y�ҽ����e��ԔuP�Z��:� � P���
7c	���hﾐ��D��>AT��~
�r��3��Q�+���чi�^�O�lk�Ę��Y�
�I�?ݫrSSf/쥭�J
�k�n�f�P�)�!��g��igDg ��z]Y_�7I���C
7��:۟��н�o������x��n
��j��z�5]!�@?���J�TpO� �F���B�DÏ��Z�:�S\pl���y����+#u`�l�fï���L|zZx�.�*ca6dJ�_)-���ׄ_��tU�׽��=�?���%eCW�yV5��
nWN�q8��xf��-�q%����q���-oW�UK���G �@�39]�����B:�;k���o=+��l�����w����w�����L~�Jd|�c;����T�/��Wի��!zVe�L�/��t{·���Y�}T��x� ��3f�2��r*0l)]=�5s��z")Xb�&z�.[��:|a�9<WP�O���� ���jD���,;���F�)-`Ew���v�p�e���>צqV���鿖�&�S�JѤ�+oWڪ��@���ﭱ�+L�B;�.�Eѭ��#I(�?�'�F:����#M�o0/\(WV�3l����#;��e��Aq���G
��)O��Y�i�.n����!�����|����lWZ�D��z��х� ��*Fh�%ߓ��w��_�d�ty���H�:�j�6�5�]irdJ-��+�z.Z.G�����z�}�����p��[�ɦ�@n!��5n�e�����d�7ֈ`9;�ʵ
����r�'�0�}4��|�x�ꮴB_������!�W�u���5�帽Q+���Us!{�^��*&Y��b�W`�+�S'&!�%�.l�c+�`.���)]��������NӪ9H�v��n�
�j���U�Q���>ok+�~���2�'�K_@WRr�d9�MZ��h��4�	O9��_^.C���A�-w�-�p����uB-Ĵ���m�-�ff��7��2�12��Բ��8,�k��u�0�/������d5��CKs!Z*���4��};�d)�>���1�A�e����%W���Bh쭺��`�R"+{�x�nh�L���������Q��"�uF^!��cBm,[x��o@��@!�FY��&��h�Շ���i�_�uO�B����h�h^�Tt%�A�� ֕�%����	�A�,�d�x/�C�1�s��Q��I�5��-�(h�qR1^~)T�bMx��n��8nrn�������t�pk�\�PZ�Ò���
���c�=���y�	�GT	)���E�o��S���I��;� ����&+h?�l�Q+��yN�m;�ZH�O[�べ��!Q�������VJ��� >�ee��mI��Se��y��Lտ)az��Ġ�U�p�D]_��#�,R��01�sp���H�iG1��Bp�-���	���m��Ħ&Z��7^ɏ�h(�����\�q�[-�,��Y(z$�g�F�Y�GA��E�7�������%���m�:'��N����@��$�4=�\�(��c�˸A� F�sa� 嚹C�FS���M�e���,�k��U�W�<��B5_7�R�_,o��J)�t>�~T[��g<�b|���w ۪O���-o�כ����������D@���;��,��72����-�ȴ���	r%/�*Q��L���o@7%��x��($�;ʈ�u��^bDH�k�/��7��B�d���G?ݨd���#I��w?$h��ȶ��бH�H�2������`���+��#��F�i���#�Z۴=q�-qf�!!|��&E�@�iW�[u�A�g��oe��.��/��19D����\��p	���m ��$�9s2�;��t�i�6����U<���������	��'-���a|,x9���\�vݳ:�N8�Dٵ:��*&#Sf;~5@�ŝ��*�U�Y\��_�Bx�|���H��󁹗j���K����,$]B�&�jy�6�l�>78�d�ZDr+��oG%�o�����r��K��1�M��ЊJ z'zx�O����G-6��3v)$S,\V�9ځ{���5m3��m��V����`c�;�%�~�s�n�-�����{����4�4�{�B�`	}9j��o!�
k�O�l�3=����0�k���h�٘���כ�p�!��HOR�Iդ�U~��A�dg��:�7vfr���^Z�SW
�U�*X`��P/��Y	6�\�S6�Nm�
�r$3\e͘�P�䣚 ��Z�M}���	�U�s\�2�^����%C�K{&��ۖg
���iH�\0ɼ֦��M�Z9M���ΨѪ��#X��V6x�կ���H9D�{j"��}L�L��1�pE�[7l4��	���}�a�?I����YA,�<����C��S)?~����D� J�����d����O���E~�A�)Ƒ��Ka�0<�#��SsU���t2-	q{�уxom^�h�M����$;)y���;=�����Os0e"ku�w��\⩿&��F�/�y�ҟڙ�D&7; C\}�!?r��57�S�=7��!�&��R�X��dՉH8ہǲ��ߓ��2�l���WC���E*����"�R���.�)�e�f�"[ի�"Ik������bU��Գ��-(�L�3�u���嬳LҢ,�@���)ddf�oA�[�����C�T(�l�;C��ﳋA��[�o���t�d�~�5�p�$Թ�(�M�j��U����	��O�������qel\^�r��KT ���ѿқckѨ���J�>�ٝ�r6�N�]�S7�YX�8cf�(��92�"W����ş��cˮ��>;�P����$�;�;N���7ݫ����ٿǨqj�UgrU�m���P¬��[�/	�n�
P/�����d��%{��H��*��1XӇc]/n�~�P����b��ۍ�y��,P�r����_��e��B9e�#T�H�_�1����F	��X���Xf@ ~��H���@�����F��`�Ŗ�[���Ck!�g�\���+ߟ��Q�<ۋ�8QKv�c��J��$VtF�Paw���%3�Ã���So|�Q i=P׶X{ ���o�B��$��V��g��
	�56�5���qT�ݹ��F1�\< P&��|�^U>�9/6r&��L����ٍ�}|lX�HdAF��ڎ�:loPշ�tkTX�4��Bd�R�y庺8Yd�r�m����:\�0�:����ޞn:�j_\�;~�"\��\v�F��}��P$��{*��<����i���/*U��v�攉{5`�R]MڹעWikv𲖶V��x"�X`Ƈ%.��P��ô_�"��U�(�b�:�^N����Є�}4�D����^�3���b2��Ks��ӾF"��Ϛ<��Ƣ:F��Zׂ�ρ�LJ��ΫAK�q(��>c��Ţ��������U ��[o}$�^D,c�o_7X&07Y�ڟ�S�^Ċ� RV� ��w�MQm	��5�P�f����$\>��Y����Y)�a��_m%�`�+�%K2�# Qm�3��z�V�g��:�r^bŧ�6���b�'��?qC�Z_R��
Kw��Sf��}A�\����|d�~3j��O~���Wp}I2c����U.��~͑0���ﳖ�Q���+�����R��:E���}���8��4�c2-�r�~ӆ��:^eQe�4��&�f�e�j�}喙�51_����wT@�]r�M�s�>(P^F��O�����*ħ����]l�ϑ>���r���'���2���1�6T���	� 8�-;�6���A]��{�����철�dg�]W{UN745�i�l���o^?t�x,.��0�(�h���J/v��y���B��v"Mg�pc��AՅ�U���z#Ф#�^�KV�UyJ�*�C�j�NC<�j�#up���y,���|p��2L�8!���X��f�L��N)���Cs#*��V"� B��[M�wR
R�FË���S�]�[c�q"�3�xU�M.T�mC\�dm*Q0�5 �"c%Eׁ]֜|���a�w�caס\�KT�v:��^�I�V�di��T^����7�]'��I<��W�4Ⱦ���湕�������tr�fr����S��ȡt
��d[�
�A��0��WB��]�&�h��?~��7M�Z޶f����T����U�sW0��
BZ�j����ʧ|�����\����A�eW�Bvo7�I����Դ����cP�
�r��O��p\>�����h�D�:\��>��NQq�aAx֏^����\pBzI
��L���\Z����z�z�d�x��ވ��:	�'��o�(SԤ&�����{L�"�:��0��'���>�%���l)bi��Ъ�^������d��*o��=t������~mkW�UT�~e���~X����:��g`����SA���
o/�.�#����	�3y��bj���
�`Y��L��î�4�~e�U����Y�U�3̶v-q�iq�C
=!O~��ղb�mEא�j���(����j�����_��n�
ubxV��+om:�D��%6��b��a�XfN_��GXO6�6�u_�||�I��g��*����<��^u?6�W������}'-�%��m���%x�be�"NK{N	��r�E6!�2�� �K�A����̈́�S���Rwg��ҝoy�6�dJ�]��;���Fi�C��ÅVN���i��M���ŏ]4x��:�R���h˖L����:+�䈁n~
��m�Epj�JJܣ2��[�t�g��V+	,�*�N�����_�����QI��RA�bevo��E�" ��$�*E.�w�ļh�,tD��Wɓ~_�d���}t"$����B�vL�H.��	ӇC>��]U�J7�`�T��f-g�ɂ�������v@�?Qlh��p�8a��H�ZH[i��z�g�)�Ȱ��8��f���t�]�(�x,��`�/�lL����o7%�̂i^��48�W���{����`���To� ��k�V핀�el8�Rӝ��ϑJc4�$^�zSp�R{���� P�ʐ�\R��=8)��Y���o!pV϶_��!%��zAK����"�:�1�{�8Eբ9�!J���(��8=�wlJ�)��a�����n%�R�ijt�)�O�!$��T�E�K���P�2�7. ,D�:�N�����ƣ�4���y�*���D�8�F�xY-H�PM\�L;ǖݕn�rz�*�7¹�\�������@/��[�����^b$�?�ns�&����]K�hײ�����Խ��@:�����$�;��YF�IefSq;�����A=�0�v�QPKyS#l@�?����D\4�U\@�f�aV�%{����V�&���V���C�n�b�M�\"��߯�EZ)�_����~���r����
	�l����D5݈I(��L_�����A�y#哛MS̬�5�ڸL�V��#�>c��<ϖ'���z�z��ܲ�HY��a٪A<#C��\pQĄ�Z����,����O��C�_�d]uS�0��i�ٓ���.0�=��4j��l�5P <L]�Bs�x�=줜 M�y[���A���*��A���6��ė�_���*
�o�|+���/b������
1f3�m�	�0��. �����Q��Bx�Ld5H�-P��=�ŉ�R�r?}7ٴ�O�x���(���zrsj_�)�T