-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
OAtnrywLBJX3FD1Dlu0C3VQwNVOOxh9NAp0cAggWtX7wY5G0u+2jCKlS1fR5MTljvegWY+eEkQ4h
x/Q9ElP69tPpxoYYEW5AttbQqxR7InfjS2YTj9POvpgXKalRiEoDmUAWtfzl0ytsF6B6jagO9K7Z
Fh8VYwEYYTVPw31yG0BKciKVfiXUQ6BMKe5Q//ZSDL5b1m0VSMp+xm8KW45GW7zaOsgrybU5kty8
SQlYcWphhhGjk1A9cOIfHp6vsjqeaImta4vqJHHwup5u2WaWwo1qRtY0fU51LuEJ5CHBYK/W93SY
wA54CBiF27xlfh5ZM3xDl+nWpSQj5Axj+U38tQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6368)
`protect data_block
6+KJGvSFriX2pM1KrykuKfsz0Z4UUDGrYqMejLn0ES5cTnn2mUML8UUu0ZsYjY5Ul3pK8g0bJk96
zfoa1JwohFThny273t0cW/3duhhajg2V+gId9DJZqiF3Is51fl4w9JhH4IKTL1ZBT/Cpuv8ClHi+
7HQF8jVHTTHbQVjcETttthD+1e3gSSUUmoJs641ZIwqxTcliIGdZrt/vuvKWgJi0Xjj26DobQtp/
VmfEipAe9PSoPQNtq/6Ith+2p5N2BO5EqPPaI2ZA/M39dEHjwVnYgNO0IDKFK55kzHSrpi2H5w6V
RVXG6wIGqXWNW9Apku4nirqUcLkaJOW9pXKIy4yLvowHVTbnXCJvhLEPb/uwKDL7KXWhkoZD88FE
AgORvfcYHrfavhha5jq3mH/CLFN4c5kl57OxSQ0U9EBRaBAnUDcgYynIyXoh/HUegm7UfYutN/dH
v6fb7QnQSdvAWXOVbiWV4neXq0DYmlYxaUm+G5gIfO+ZmQ5A+cpoGJOX/qObs5jrxWo6OfmybRgZ
C8Y3JF0bei7AFx2mv7JevaSH1LDCC5iCQt/klH8PcHZwHWtlDepXdJmZw4KBGiJzEmgZxULSsJCV
u55t4RZlCqfDmxLut3UJiA9h7GUA3CubRuG2boHBB31TBnDU73FTKqq0IKef5M+Eg0XVF1fIMnaM
A5HmRkOy9mOCEKmbkel4/mNS2c4P49x8+14Rh+6kv5PoEzBv56JD3XjOtX0eo+1wBCvsLzwrmRXi
nrGXMocUMZ4Ol8Vo2nyjy8/mDeFRbCPesIxFq88JfvWnVXOjnU6eBEuju0ojMeBYQZ8NEEIIrGjP
dbMuyck8ywvGpcPynwZOMqNqMcYE2+1pHoAneKKscN7votYdwGNfpSmDbfK6gtZTkpCuD6ygrMDe
5vXbdJ04OzbksCbzqIc4EJTX8BwU9gYU2O6gR1Q5cmVrJ7LWm58LhxAqaueaJg2hTDunQf1+YK6v
/EDcp6V8/iBQBGT9GB0IrRxQ2fOR2gRvO3xOZoe6btZJOWF/2yhM4b/8gvHPItziCNMjkKwqEvd3
wu1y2gAk+KLPtUfL02n7phQCa9okEj5BcNYmJnyAuOVXk+EpUCaEaUvq3LiQXIUPoM7NUH7IutAn
EKoBV5SgIFt+2wQLXp/Z1dVa29Fk6vfZJ+KFEO0M2b44ooj7OPEAoDzFysRLegMINrAa8gUXIR8x
kd5KoyTd952X8JEsIOJEmERBP2arrlyH33kFJKiB/nwq74yUESSXlKyzOIB6m4T78Mp3JWt+N8Vs
bkL0WOWGmuCQccE4Q3MfX4t1gw016ihgJdUyOARE6fIlouFXYBSRPovZW+GewPPoXdJgK54fp6Kt
z/qfMWJMfg3AvLOE0XSoz+otAmMJofgYyytLimYtd1FmMipWP29BEfGZqmTViBRn/rSMkPvwlit8
OFs5F8hlvTOpMZ/jMeu3Vr1vgx9HTv57A4bqhSvsxtOKTLddCXaspxwI+KCSWaiD0w6DRSwU3257
pIrpya1coyEh2oceH5fpIsToHXG8uggvAAY7KETltmkm7dLRzIIjqNWKtIkBnAi4isXC3blmxf52
MT9CWRIWe4VCbK3envky01PUPeosoqP7O+1D5EdD4zKOBiBrVZz/1VPiynif/vPC6bsJ4eMJ1LPq
gk/7P1Ip6XXqkV+ylbDGcYQNmglJ5XEFKDxcMW/Dqo66lLJ7pQOlGBc1bZtGcoEeGl8H/c8a0cZ0
/hCMJcConFbgy5vXwi/GbIQlNiFjQHYTzp91/pUXuIKtNWHHSQynrDRFSCgxdYqDMN8fcDQX6WLb
DDyznYv31Gqy7OaAO/7NbrHyQllej+pQjhXnut6c9+rh3OEd9ZM/xpeG2imONIgLF+bPTyjA7peV
9DxmcP1uaSzO7CfcxPjkQT9Nc+BHUQXGqW3ogRfykQZNQjQh7XYKtHVOQY2cWNMx0hlRfjTeSRTH
9d7wtiv49yvqd0bx4pO360USN2YmJSbH3q9lSKWjKirUluqjyltBVkyqaXINFVpX07lHF3tRtckU
7pCS+PRn2zkc+9w+SOhOC97p34X4S8k+dpzxaQhNHVeLyto54I1p61jOYRjhJ68jhqchfq6rkCVn
HeQ2zzeGZTC+OKc3uJhNmlCFLnI1jjIvM6t711JBs5u19joUccO65HDmX+rfGxhiaas6BZWj0TbY
RYLwC+Q0UdA8KI8QJZTHFiCHbIvntaFF0DA+TZKV6nJp6xt3xlenSi4yWHFWgBWzWpIPfkEw5dmg
H3o4jT6/LJmYYmxtWjwCJUzXqQpxDVQlxYO0KBQkEVc8oWrVFukv93klkPQMqBno0b1yQyXh5ytc
um2UaQFRR+lO7g99l9+57/U24N997ENOhlmxlK54HolSGeVWmDjvKH+U43iyKv/ZlPo/DBh5JFkn
vRCXr8W3jSjQpMCHsvP/D4MKEqQ7FUxs1xyzhPZ/ajBx24238d3pMQvWg3KxdBCVhEdx9KG1lhGW
pZK6GfXdUVKC2zn2tsRJjrQjNsx9BSFnN4knBFqpDlg6JzhdMrRdKwOHkozfcT3E0RdYWEqcCZnM
Wwt+aCYZB7hj3LSgH5SfnxFYELacAuPwG7Qo657M7vdMjOtEs9aYtX5S5KMl6bHj8WlPx/smZwmi
g1qVJGxN752rzAM/FbOyawMSBrXkKKzkUjmyKVhbU3PNoVBKuylMfv9QCmsVoWG940lsUMiRKYhr
QQlysGoIYyi9pv4nI0UbgqLmUQPw5k6QNXD8zWJSBBpFNY7OGmGROeF/k9SL48MYi1LkMaJNpAyj
NfbH7aXfxDmTwEGfZSlzHJZbAd7yZdhykN0F77EZZuWS5mcMcFPzNi48kKgVZWoQJdxo0QV8Stub
UIIh57nCGVPG2gGQzp0Wrms6JkaiZ7MUCoJltC1W6nxxG0fH/ub+3OOyR5JQbLj2O1Vysd1Vyutt
aZpozf88NhzBtZ5NxAppKq91Fai/Ig6h9Buf5aXBOPKUlCestwPFbzIGMRBwNFGTzouMCMxPwK7i
ses10fN17WdzAAPZLzy6fQoPUjduM2NRiuvHhc4pBjM/A93O2l9tYKjvSFphC9qVIVA6+Q3Fo7+n
Oy6L2uMh/bhyo09uUJelSk/rwPTDNoFQ4tJDUNFfMUaI6S2hR5MhbRHzbkL/NdfqEbkC0GzMeB4a
TfIfT6ZJIQOOMXVB2ZXawvHhAnvDTyOF1GYzLF08g3EvblsARmCTlY3cCpGKB5ke7X+iQF9nvmti
e0Q1M7cOB7xkBiEoIxAXcEq/mKD77Z7QuiALJ2a6/Iq97cerbE4dWTDA5Jd+9ZCQUHCsJvcdlf2a
m4ik9KZgv++IagodN2YORBafS5B7t6VDThgB/H1pkhAB7L4jDwYSCx+VzgyTVcCkqutof9q0EbBz
L0TcXocZKC0aOoG/08qTcdFadpZHo3axbMupPMZZlb8GJRyDNDWaJE0zQjX2wpjw6bfI94NV6D1K
UTM3b7qpjM/MbvfhJGGg5/2UPSaE6rhcLvDKW0C/GtkkFH2OwZ/COFIgeMLd6wKvasCS2T+qgi5U
ShOaFeDYgLAxhuAWzI3xZ3r1Fp3tOg/ut4zLR0ET3k4+/ll0S3Sn4VGUcYDLWQGlmsfgGv5yHqzt
e3i28N9sqeBO5zPuIiG72VPbtLHZfW1173SsaOGlSc5mYLCyMevEOAIayta/hv6H1lrfT148h5H/
N+OuuHm7Hfu6t+tcZtmo+M7JMnBuRmQyWJswMOaRihNo/gnb2CywApyvcYSWYO6FKbPrIzhYpeT8
NxJhlQJ5G9TEGmlXd0cLfEZMsY/YeJ8beyT9lYF0sDCmdjvubB9I0j1KzjHGyS01QpCAXWVHoB3V
AcFmEFsBCPcqOM680JSfww18KAXzdN4psU1R+IzQS0/ouApN1+WmoJdeWzexxN3o3ynM3jr7HuUf
e+eDi1Jko0aF0Pw7cv4tJn5nYk4G69a1bYmsEri5mpfVHNd/hREXGshFO/f18fzh/qq6CFUomG6B
BgvRR9MN6Lj698JgY3mXS4VGMfFNe3GCinnETOn8KxVAGzwoZR7VgB9h5EpcwEnzgABDaCNjYo2y
QQlisJQWaMrMpejcHncZgMX9feXCa4OVpo8GTC45ax3KdgLXazbQ+qm6NOF1d0vggiYmvBHYAz78
T5Y+zg+cz3h2nTanxdPrvWnnehAojAnG/p1jesTQRCHgsdM/NZ9hl7fLRGy3hIykphc9xvrkaXEV
eY8BWzDsQq1hzxsOWke/ZlkyFOZK/ZreRNZoNeEgGc4DfjMTVDhiTBHdgDuQAddwP9sm3NEuu215
yEAAhNrYnlJK1Y/PdnlX3BAC0fwzU8iWdjf8J6H1FPCOPEepe5Voox98Zj/7TRFr4BGoCcBF/B8U
sEysQIbToI09H0j7pxPjO3JsPm4n9ZjjVaDeTYOy+SLeXZdo9PpheXBeOrhhXTl4NR2GfUXxY8OH
mNk22BYRYDERw90Ae+AT1lmd4Ty36OdUbrI7INIltgBtidSUpZ65vGsWxZwBUqn0XaLK+K6ga4Cp
Qqd4IiuBALzUkrMSuUbHbqtlOMdsjKhNLT4+mXSvHcd7tf2jpf9sjFUmkbyXPIxBLH2sEaOxORlm
NlYtCF1BGkH3l7qgtpbRAFu4ZnP7ilqlUURuGFoAQ+VihohS9sDw2VutfEiCjeFxmgJvOsOuAWkV
m02wc7HX7x1fPbd/eukLh9YBNY3h5wY7ChKHRSl6ZZ7DDk4zKuLJoZWrfRhjKIyz4iXaZJS4C/rC
/TcPYB479znvOrY5giJ/a+UwrCDdnHUDI+ZQUjEq8pHgdPB49Rnj1lpjbnu05nYovq+16Kq485uI
YhHyamIdU2oJFFGsxsarNxjLKznkXGI6R6rBTsGiB1ih3ilsqmiQ8uniKTrj4zpLyMZqyVOjenui
iJBe63Etf2EuXIUW0gaZMq5YOwXRrxesLjAh5r/pYTZlxN30XYrG6o1F2e2P5BiWIOI58KCvTw1r
1g6wQnFPJBjatk9FKEnWknnLDmdru1ZLKSuvz2x2hJQxFTJ6liqil5y5pJ6qF1xNMuYEJbwDVINA
hrwyPvfuI5s8s9Xous1wPDDViY7fSHkKgDeFNjwuaVvGuvXm6bCq9u95zwZw9/PYEj/42/rPgjAv
kekDs4BmkkVgLVvgStk4h1AAbaQWYu2pRVpDp97wrRh4mzy+nDQdmUi4uYJIH6+h0pLglj4PEZ4c
6vKuOBjK/CD4Q4NPl4MTd6mnYIzEotzNnfgm26rD3rSt8mIi5MOe72rJDTYtVqbDaJ7B8mW8z6bd
8vVBcIjepyP3lcVCsHqRV53lsImOneFWg/mdl5N6mhZ9exXsAhGYvjaR+uZe9Bxmmb20HyhWgltP
ShlhNh3M9J67yHI5ljO2KjZ5nT5SwxkL6eqcWmP2kB+eP377oTjpiOxFh9LFy3Hu7lzwx0hFG4qC
7I+G9KcnVCSux1svLZxQRfQHUn1+zt3qpt5Nnx7qN4Pd81+ClSn/yySOLOr4gwrO1hswoFdE9zxd
ISNyIujrgjIqxnAxSyCIbMgkCPca+4S0v05g/96bV7juwzJYJ7sOSGP8n50SOu4Y3DNPjnnaqNli
GVUBbZ4gRkjRu0beLZd67R7qjwoHRdWR/ByE6uOxbhaf+1UVIPClJ7sj+AVXhdxKnF2t2Ohyi3la
XaLFpfAVWygAd/aSBGn5sTgqvVKvgQu+n6ulD3hYkkt2MB36utxzRGIlivZsna9uPF5l59/cIYBy
onEQw72uEHo7wqO6TUqHKTbgINCgHYkon/swqSLiaU7QUigQohTtDT9JBFW4H/iuoCJ+y66ZzxQH
AqYlcK8oNxH01YBOd4FQskeNoQbTg3wgEyhJU/hlWzOo54VYn5/YGu3rZzEheKGLG5h5wHJ9SYv7
BjFd3HinjkdZh2UhkmNCdFTj0OL1B+u0V0q9LyrXMaxDpGeVOayo0f/jrlWWCWs2QN47hlsLHFgb
8FvVHNk9wjN9kcGpelEIu85M3ckpJ7KfXDVLf9qNNmsWRFsPPy8vHBq2bmRigjLB/mYq1iUZwN2E
nvuhALgFaO7RdgTkcAZOhysayUkFR2SBOTQiyHdP/hWvByzDl7HK14UkJXDxB8c4TibNzliGGCyE
DgBPNqZd7xFzVHvX5ZNlfTxisqTAA31n2Dgbcv5oGWccCLoo33EjP7q7oNS/gu99eDGbFqrZgzA/
sPWELO9qDZBL3G56zOaZsPn2g9ol1k68ofyCfX9OPU+SD1F9bDBFpWpNNkGGAx3B3YEvVtrYiFJM
BoDzrtsZXr55n0MUvsmRS8H7wBqJBddDOsPzbmNuiVzX1Jiga2/0Sr9srLm+ejRzGP2pFVUc2HII
g/ALESdHsJOv0k86DFLSTB6LKOm5hIu7fNTh0+7DQqFlA4BJEteLn5UDN+uM055zXwiuMsmQ5LnJ
AUhzu9wf97hDvYt7tngp0nHA5ccC6umt4+SX9ROirBIg9kAKEu4VJrC9K9rf29yc2CFR/v9TrWRj
kbsta00nhAPB3Ci/m4U8ANYHzhHrK1o2mV8korCb7xc2TJbMxJJjSWUBpWER/U+nEht+9JnZu+8+
FplBPB4++J+KZJl+M8Vh7Zd7akrm/HUZTavvRq8oGwPWg7Bg5yR3okk62qfZdLfkWLJX+0NYGyRr
cNb7+3hbF4oCavPcf9yKWumA8uFflAGr8jSYYjSJpAdz6wkphJLtFKStzFDaFaGV5KwMOqmz/Vbl
Y4bOn0W6N9JArBLEmDkufA1x5mnt3Bhkjt1JSfRAgugZj+x28ZQxJM7cV2GpSvhOWBUd04esYrjo
RwsoOzPLGmlnRO8VUYAVGfcT13+X8uNejAyj/EjN+O7cFGiEkqQLp0eGaXlB8m/2QOX6Y4+VOODc
kjlDll+9ZOzbYDOI/lXjrluRwTwzrC7P4vUz6W7R8AYLX74jYVZ2m5IALIU35hWOut4/IipjNAkJ
a8LNxpVpAZNtiob3PKjYfPSxql3iB3c3co5vswvMp0MNgVaJQfxjefOYOrUwHyqb0tfShmVLjl1v
fmJHkqrnWwf4oMrAt/LD/zEZgVLNkmHXGuK7lqmWpPHVk8xy15CDkETPiOqNKNHki72PktBo/OIn
8jK5DazzcfC/TjhSqfW58WNP05X5/5OPw/l4ZzxWBhr3nOuSDAbOGQ9uDuMxboPeY/UZqefbeJHS
Arxsz9WB0oTmNA6w2KW6YZEI1sISmWSV9t67IYKpgVamf+iVJTxHyIm0iMKMz7U33sfM6diidx0N
2XYCDzycBIvXpBX1SYb/XI5jZU/8XUeVIPEqkFUq+lg54Uq4Kt1aQBo3WV8mFFLQJdquMCORcJr6
qX5dOs77wzfUoEWeidbGprHOjV1PliZzG2vEhKtH34Wkv+1B1hbbmhUz3WKcGW36gFfk63rF2cZC
c6tCc9IumBWKpFHanKfnQ9WGt5YvWonY8voNkdmfndwYgSld9LZbmZq6lNBVIHPMk+fFQ5e65Zr3
dCfQ963PiBG2Wxdu8UMmYlOVY7sXmGE9/C09gpY4QUYuPrqiiGtdI1fqRgGBRRhXWw6UDYihb15K
6k6OWjuMXdYqJV/yB9BD4nxnSjWp4tiK79/RGXsm6tB0G8NCv+t7HDz5KjBYLLQT2QpwtgqTjog4
AaaLg+GYG2rVM4jujQCJv55Y8JeWZzAdsoH0SxYw33kr+flX6FJzh5g+tFOQqu1ac4I/O0W1fKgR
c19Zg0lv7Z8g163q6BdSRKVJrGTEQtAV7WE/n80XQxTSYI81xhA7s1iuBQz4U7h5D481iKnSomaF
BKmeHJjIfgDptI2b6b6FOLCGHzNSif45izz00I4NUlhbwHeRK+aIATisJgehBv9mFxSRtX9/BJsm
EJSyLYYf9tdtdGSh3GqFWzddgvNxgnZ/xw8IUhKQRIOlCQOl85tFqDbaFY2FgM6kaAwb0q9bAtY3
WlC6/GKqB/nIJsLgwiQZ4OL9KZ0lg9Wd3RibryBK88Zbr22NtBOb/HT5YUq9RTZx1TnsRMNSQGl/
UwecwcLCv1raHcCNnzbFdwFOu96ydbLAf8KlSkwb5FAFinaG5yRmqthfUuaqLiOFIpOWYBHraUWo
up4EmkGbMDmW/q8rnecT2aThi0Ac8mCH8DBA4I92F2pfyBDLvi5m3j1yWHQypYJ6GPCNSOO0YRvx
ZCFIcG/O6pf5NBWaUaBBc4lOJBW53s+KTSlYpdlbTHF7wrxTP2ySl/pJSsV2SPuqTD/VlSlNuiQJ
0dDB3q0XbrcTDIJbX4bqpGS7JJo+soz6aAbEse3vG+yp+eGOS2E7VktzBrYLEDep1dat8MQL3Nzo
xxvGgCA3LTs9t1GcuqIhWIB9Jq3PC+sGPjy1mnAaUA4JNzDSdQVmRQzS0TyKA0UohGseaeh2pN1n
ZRnEJ5T8YqIn9x05l4UY8ZEMEtg6gXGZcfhOhzo3vWoyuUJsut2IPbM=
`protect end_protected
