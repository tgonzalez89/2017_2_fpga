-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
rzqjxSmpFNaKeKRMqmXT6RM9n2NHUlqCCiruFSI7ZRniex1WuMaYsu0K6xhU/yPJxAoDY1cAK6mx
o0UH3NipmdgDe2bSnxoP0lAaDB9B2DIBECJEaXpUlv/Jwpitb/KBPOm6qsr7m3W2ER1bsWhQulAD
an60VzpUMslrUYA/+rWGV6oXL1Qk/hVwkTkSnUfEGVWQXc4I0JOxFvLgFZtSXbSzd9QBL1GFdtmo
+jlQvYrXFyHDBqDPr1ios2HqbmghfKSPWffXQkkep/03c2/aggDPgtJO3F4W38dL3sO164XmeOLt
yP9NrbmpRiFWdhGV0G3ukJmAx5FN8Hn/i5izTA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4832)
`protect data_block
226gdwiw2qxN0AiC8kLtciLM/ld5456SLOpbEE1QotFGpNviBRYAO48R7UmR3UBpwGAqHJWDaxzv
6oWheiqWwy3HwLw0aB5Fm7AMV83SkqJ34hWAuNdDMpA+X2N8KcHUeHuFzzaDVZU4WsqxHAr0aGN7
mudt9xGcqg+NsKagSCpjFRqImkfIRDhvAmLpzNif9ez52Gkqvk/EgKWrbRCmqSCrCbV3WTE5dBFX
jVVH9WxHFVcdjsuCzTdxnBLXMkmkJd6kIW+SQDyDIveQ3DsSpKI2r2IykhyLxDiOHBAQ8rTKxvJq
Mig+7j8nnlrIZhdsQoZ0cN5C+0C2QxzxNJqW0hy4nEkDvP13rWM7FboJFXyUm2mOrCEhM9E1MBsj
H36qekCxiEAU4d6TqZYALEKdzrN4x72w2uJRqNZ7ZaMSBjT0PEpf9FiHeUeA2RJ0qDXD2tjbohaL
ezHb0MK/yRYffkMLxwJv9rJvXtOEH2HNwF8c5OLmDDpsR2Mbvq+/JJD9Ie0MJGx82pbla8MEnT56
38ybQQ/ra1cnc+9zqXB5yLDWdpPiYqyOCGAIm6eOBJRgPdQ+tgr20FsMtS3WBYGBJ3CGbxIfeZaO
FGHKp/DbJZ3vPu0hozcTs7GT22150HqDwWeQqXMQmRa2uPD8CdFOr6d+0CgTdyKn2pJPBSDt5OEf
1NyT6kdKn83XDgYQRCoF0mr30yO6EgQ4LvkfUITcYZ0V0EGANcLidp/3wg4RhOMMiXDbnOzLRJMm
EQi7MsLJglVfvyPuQppbWITsxHUTrTNrNe9a7O5eu2LvPskWFstD7nOqmBVkthkLzbG9owDabP60
hiCvfp3zevq+gFk2qlXuVMl1KLCe9nBoeFWY3c9/6hjiapqCg3vJQTvIhMJLL+BuZ90KzYL//DOd
llxqOQvoxhKbLUfStUxE2mngrP0PfDdMpGWF9Ze+gcsrqOBEH4HDGrgZyZCm8Z0udM6xO29Ismsp
Xy4x5fDAbqXBycwy6TUI+GKwSaxkaJlBDBy19juXtNRS5MOVLCelaVk4DYlMJsQpj5CQOtMSvSYs
JdxMmYrikrpCsSYfSA7QU7L0BPAybihCgpuaMnmAS/VzA5AOROdT3t7RZVNbfch6mCHfsWazabsD
hDG17XMcF/l+QkMui4Mei+4CsA9knOVI88J/60nYYqjK9+ZvvPmXHq6G2wGQwqD5JDWIuu8p6VGG
ETblffPBOiLTOLrmYNu878ttTbi6rFf0L58UAWM94FtKE0IJrIefYcKdIFOgEjlpLEvtFqk7zDLy
nqEI5Zs65AanJvKJW2gQCg9MqawYzSjWUPy5ytdX9q96rO2N+A/bq7TZ97gctAVqgC7oJc8ayNKq
LmXfILhOIjYjw3tqI9jSX+ogjcfSRi6ADPPGAWw6Ydgh2Iv12Dk9KVBWKvU80FHNvxtJ7TQl1Zau
pqoSTyS3Q5y3Xk+zUxTolIS7Z7MEFkLCbQRKRoM9P15oZUsW4whb/uH2qd3jqPtrS1i/zu2l7ze9
PXh2VG09zFhZ3+0JAb+ObU/7DnKKH0S+gO0uJZlxyn20In9l4TOIcy3jJ6914G075/BPEjjG7isW
pgyyaiDH0hk91qwCIJD/ce0XriPO0kgBrnwvRACjDPATC4DYvL/G2t8n9QRGJgfK4m0UKTGcGwFx
28mfxOSjuN5fi4U4H83ZNCFdG6OwyujkT5FN4S+ztXsB0vfq++jp2Y8KZOnKuigkxexauysCYx2e
YlQ+Q/agWSvJyd4Kj3KCi7sAXDZXYB7ehM4XVkLZkJN+doMlEU6mQTRHL2lXwHenhf6ZeQtCSMm8
LUZRgrT5h++/6RKPLrl4ooHurrNJaKSDH6RLDKK1sfbeW/OoV7b4WqCO7Je91mJF31fz7h3juHOn
nEzMa9kASivejxYHGrbOKX7tIrlGxG25bDLXS3505hqo7J7XcS4Xb7ltg0r1kHmEquS9HCuf2sb1
umwqu9W6Mx74QJ1sYuNu9jKjRcwtj/iwUgR70Gvn3PDeb61vzaQY7Pm5LQHnUwz7BP+i4EGzF/Zf
5PL0GCpHidgunRtEQzHLJVlZp1OwsJHr3i88MQhYBV++BHsVUTp67qIAZLmGtGPdgK0eFQtH7xRn
vmkQX9ZdPoAIK4m9ZYdGZTG3HfvQoQZTQWosb+dsAnjre9yLhjrVcGFPAIbI8oqCRNq1TNER0v8T
5U7KKm2uBYmk1SmbP/oCuqE2R33G3xq/D7dlua7y4MgY9HhffiqknCFsh4AJTGVecPJMWGnWokdM
UWj3umrmRacT9aW4JXRhGO3tURzh/+CPBKxHbhCMGzddxJMRMaezVNm3NLiczfEd/eUBVBHgJysV
vSoLmBWOlFMIPAVd6xV8vL8XrC0XKMgsm4ZA3kSA1w9JKuo+So1F0GiEAzHb7g06CHng/U2oc0ns
XDPKRlnxyjuHB6XbnnP5izK1x6FZHMgFSJfsa65HvOX0B02+fyt65V4A4mj+UkwzfiFW5eSDdwTV
7Dj99bEl3+vtoZZzx03d/8bbqW/Ry5TIBpzDiXaZ1+yWXjqMuE8HxqiJ/RJL0mRaHYeT855zfiwC
4mKGdFGll8FR0ZgtSDj8FfV4FD1Mmb4iL361j0T07cTUq9EaEGeIP+29EIYB9gup8dUOd7j5ejkn
bzUUEt1wuXh1zceKO4OmqHpKJVQqRQ6MoeLJ+tg6Z46O5oERQElk7NipED/OXe7Dk6+Pgy3XL9OG
f6oTZkk8lQfrKhLG+gBd6b10NXOApLDOxbw3Cof562oRuvS/92YjoAsP9MARjKsJFZPu1tvFvxXL
wZl5pie0NrYuQw9NpBVLyWlBGFqX9uazQ5Ezk0xfPq9GXZvbxPKAJh8OaKPyasSdDcl1mIzboFn6
fVRkdYT7yuR8+SL4VQu/Q4Wzt1C8ir4KLVp0pxs5gSEFg+QmbaCBLubohWF/0VT6YuJz+QtamS1H
mvxTqOXbkDQmXMjSyEYUOaS5X3PSMr2Pj2EWfOvQfNIPoklv10qMYbVMgs/XknT5GtHcTwaSCTx9
u8A6gZ+ncQxuGfLIgE17Y7qs84/+/KiciWkevRMEgdYTXbyigrhuXTtX49sOErhXxKMzP8YdZr+C
mSewOIRe2sc2Mu8g6j0Lh0Lg2VT6CW0v5VfnKjW6TLLThdfgsqR2ok2wUJwAuKYoaO90lYCQZMtj
2n69yO8wbHj8DWs2Hr8DavHtQQwdPxa7CycSFRTOPxj+0hf70iyl4G18qhu2dtu9wmhKNBRb+1UH
PVWkmQVX0S5gm8mzxevjXUzaQ6NFi3PnvYxpTF824a7rnyMPOrwhIM4ohpAArK6Zm9BwZ8UeYViu
phw+Y3p7DmWgSGegxdQZhVzVEA7nvIzn/0/MRw8dgP27ewsnr0jTLguGoB7JqbY62tcBWxAWPcrg
sAjx0LNm1JExt5zdXNN8a4X2WNW3jFVyzV8vFH9g4T0KIVQlHh7vftwxtsthf4IIwXnT+N1tv5Yz
jooU3ooNQaz1ospMjNZ2U893P9dAu/2jfIbk8mkrPqtyjQX/Z2UNbG/11Zrxs91WUsj5ivmjgbOP
eG45uFrhe1v6l36ITlUslRDlRRtFIvjXQeo9uuFUHvghxwZKV20IcmsZK4cjF58euBcu1S+u0vcG
geXm1h58Mt92u6g/wwuUqC2mIfm67qQWRTT6HpdV9nIdzBA4rKeVohBCX7qglCyzDxJ/ib5icpa6
G2wqc5lGFyz70CKh07EQOkIRyIZKrFkyE1Tz49Nlu5DYSQ7BVRijN8POjENolx8iKoptYAvui77f
/ZZGh/iwz4IyE8xLQEsuu/tFoLrWk3sT0TlZ9kVDERXGKx+fwTF51qswZb70ZtO8H1XWBvgDkK/a
zv8+G4GOfvVj00WDFL44AN+2OdgAAkLxPW82+oDkyFqRmnM8oZpNwP/TIjglSykG885AlGYSnLag
5HdHSHqDGKbsnJTZZD3ZrnRBfpYgIlPrcH2GzjzQSuTlnlNN6QYoXQj+cGsEVpU6zZRiA7J7SWCN
hfg84XGbGt//bmdwajyKCLBlvUTdqzqtXd5rPyJezvHswmBwjZiIztr7xEZjYbqkHIRD5KJsyelw
HckikA0N2CY1BQVZExxy4ZAWgdewU96Fkb6F4ImpY5ggJmA87xAl654s6Jj7vJLVeIVUcH/23T4Z
ENmgv1SwigUbV49cLgtO6jt+2KvGVYjBn2GafmAoPbbH699gXAT6RcCB+T0pV9dJR2Fjc/KY5Ju4
l5jpmbbZQSWC5YEAqWKPIlwBsjqSCycu3sM5chqqhrt3Z+Zibs4J6nnJrPy4D0aM6NojD2KDRCkI
LGkF8lVOZ1PjGyH/HAerQDQ9lkv/lQXabYdJp+APE/ZAre6jvfNZ6kr+bwTDHvxF2uQIhz/0mk75
naQk8BZAgGNLaArbADQRC/8I9D+Sw+Poi6W8nluorrecnkzGGIRtZ+oykvCJTqeTkykkUBkciiqj
p5+AcYFlsrfcSROqfrp2BvWiRGnhpG5HR4xoZ6NfXrnYoctLi78drzCN4X+MiGb7/SXFppTxaa6v
j2lvg3RibJx8Ifrp4etyrD8s1bKkrHnPa+uKI79igCWSZmGfUk6q7QcYxSUnMpN9rdYBmWXZ4QnE
YzMJuR+uT1AnT+0RlAv6tLNpoMFxv5tDzKOQPOqyCxESuy1wYzp7cX0oNSLfyjT0RRJgyTzWogh6
7mChK0rGmWbPRJed7j/L/V8geTkq6l51OzC8gLxjVYO9Sz6Xy2Wv/ONq2xttL5bK7lkyIVjqoFz6
xgdF1adEJAE8hzHNNs/MsVFqY3CmFFBA62ZsJglAFbU0k9u1BPlezptOyv9fWRHAWTHkFTHuEEbb
sW7qujl7BHjHlUxPYnGyNYC1UaU00yTIpWzzU1tr3UI/IVfKCA5ZZC9Kmtol5kwrJkgZ/EjqAA7q
yFtLMachC5WJfpLMtf5x/6PEwQONiWGI3tlaVspoYmNi5lul6KWVJGDa2INOrQoVN2Uz/umf/Poz
ti7p3zNXg6XSmMelprabERp0bfDF8kyQkPB6GB437ae/sL85Jy2jZtUhjoHtjekV35Rqg/IDRUtP
resj7xQ60MDHskBV2dXMQE0mRFsz9KIB93f209+YQp8BD+1LD66x9Gqql8ORNbNlPreyJkBiXLom
yt6CCWoU+dSZwZJP1K21oxeNA2ST2iINj46EdDTxSAw3a5Iv9JOKi3T3N0gtYNYY69GHBr6NWJWr
7Tjll7dQz384w249eazSKn63tuzE7AAhD/lDWqMvgGfJArYUEVxL9/EHNQfroYRwxypGWWNqFY3Z
Pg8fy4LeYgSZqvKXwgcaY/p9gMRE379fqLXSrA4d4qgQc4KveB8U7doFOTOnUhWKEgN8ZAUEl6RY
BT8ZR9Re1Ci2ahGzWDCVgM4Vm4VjDKhMuu7Jc7PIHJJ4kH2BgXec0nbeKJCxIma9gbgpLRLiGvB9
8s4SZkw9vLYa9fK5zxHWhh3M+1JVMZXcqOYMcq5siIkz++nggh6rWgpPlE614zHpBcWngPk4XGu8
w/aPBGCQM4jn0kTObYtmK4MvP96wHC4vlBWw44T58+Aezee3orHU4qV+coM60sHGH8ss5n/P2EnQ
D/nqHvDx1XUU6rJSNGeU1g0oaWY60yhlGbHjxY/t4t4OdIXotTDEOpCz7alEdCTkYlAaY3ATTGk+
W8KODJHhKH7kk4iwl+Aq6bpeOfDPAC7kv9MdeRekKTD+LDK4ks3eAMBswwsinJiQzcbe4VAlmn/O
6pM7vE4UR2e4ySHdqaxyELw7N3KThcjJZiFHUIGF0hBV5lyZOZ3DiMrlDOGp1I9hg+HvkyB/FYYe
wc6GHYFeeItUd0/5mKJvXVsBlb6ybo4BKhE19eDNy1m/7lwfpITovinPB+Mj1YJF0D/OZsAbtMN+
TPZOZG0c++UrNVFyjEM6kJ9OR6bXccrxSESLZLt6p5rQqMLnrAeavCzA34/fV5sWLYETvE6Off7i
EaQp43XzqS/jzGP7qf427ZJbnta65lAXkE2vF2GxugEibsl2mkJWaytpqqDNF76oZxm4j4ft2Mfe
hjg8E3jmTWcFPDnW4xTwSDFs8fet7DYxLmxPdOo+LPqjGhLH1cY3Qm8yRoR108GWTQrpNDNaOBbB
ha9KvYiBe6cW1EagiSSLcjCrc2Bj9i07g2h1WjNgfnYGMiwa5l0lDyHtnQCytzG5U6mlC4LvkZCn
n72QltFJ4dWWG1e1z0xzfKRevP1+FebF9BxDP86N5uezcT1Nz3NfhZApD0/hUyzB4h3zDSHYE7ZX
1aXV8KlCpeODnIpCzfH71aScjX1j3byT6E7gM/TWgDK2aNfhWnritoFiMJVi05a8NUYcXdt2xwVO
m/ooLJM/KuUd2fl//cu/uM2xhraNhYJwPOsmzoNNO5rcjUAY/q9taCbT+Fc=
`protect end_protected
