��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR�G��W������W�l�'�h���Rt^�(�F~��@ĺ$�ŲY����sv��(�{���J�x̝�y2566g��o}���z�%��dX��,��c�|�����y��g�mG�����]`��f3�4��8���R�@x�̶-�7��!(L5��`3�~iw��>�J�0���"�n����\q����$��z�@=P���56��tXx��z�(�����d�FF6��!�́d�):�9����_��u_ݓo~@��$#|�3�RSig��Ƥݸ��z�M�1�XW���l��.�J<B�����sI�S���l�x��D��i��P@����:�[V���J�+<�e&ڱ���'�{� ��-���$$R�s��d	�6]�}7�/ l�3��h6�1��f6������l����W�=5�X�`��{����~�_���K�Nзk,��1�	-��!��+�����0�ZG�9�P��야�C����0^��N4�ǜ,��8���EE擟�e��C�L�����T&� sZ���y⸶(�rL(޺�#^v_h�W�p@��BL�����K�qڀ�7�z���3�c���g
�Ӧͦj���TLL�a�Ũ�Wq������4�7K�w[=���)�y�{��uڽǰ}��Vڅ�����J��H#���Sz��濣Pe�(��A�߈�i���VY�]��2_�HOk��a�ȶH7��L�E��8ٴ�����6^mc�c�\���v���H2�֫F>��㰹�hq�0"�bκo�
L?Ɇ��n�r5��[��W�Q
GҜ*����O��i7
�;����v�̭�o;�Z=�AxZ:�淜ι)� i�J��)?�����ɮ�s�9/�՞��>�3,@�2���N�t����P��dm���u�dEV>���3A�v9�,��	�l����7�ۧx����
M��`����Y��lqɶ0,D�T�V�U���Zl��V�L�,EZ�V́1_����H��Hy�ꬽ�_�p��Ôʜ��_�g����o�
W��ͣX	����.�!�4]ք>�:�M����ѫr�P�C$�,Z��o���,c�5>/�4�Çq|�+kѲ��}��+?2#$ٴ�s��OO�@ʜBU$�I��UqN,��sd�v�ïP���޾��*�_1&+���ݦȁg|����	�"���Wl���Wߖ;�en��� ��1|B�H�`pv�B#!.�UbCk_���eL+���Rn�+�0���O������w��W�����W�(ĘUeؒ�|2|>|�,��pr���RO>�F._�e���
Ie�U5N�.���%�@Z�m�^����˞q��DIPҟ:,���c����E����Y@�{Q����fȖ�������}��ˉ*+}t�5򍧉��
�l�%��ݖ�Q���sЇ롰�d�O��釭*�Hڪ%�K�0K�g���unZ�pc�sS����5��Z�}�Y�,���v���	�9&�f膖#���iTԖջ ��0H�	{x�Qi���s��ю�Ջ-޹�O����d�U��J)�`�5�fͻ�=��\O�(L�<��f��֮��ʿ�+F*>���4J���{�\r��j,�F`��c��0v�F_,��;Y��,��'���F���)�-h�B��xx����һ�>I2�?q\���Z��_υ�D����h��:Hk�*��7��%I<��wd�	'&���Rk,�ޝGJV`s�r��Y(=�!���^����Z��=����������"d�
�̝$�Jc������c!'�t.��	B*g\� \>|��}�: �̷����C�:�N�L�98}q�����Fa����;m��z���7�{��"�#�v�>]7�_+sH�yu�\(����U.��,��Ĕ��[�Ct��7Z(�����~X�Y�-Xs�&I�z�hC.u�1m��H�+���z(��=t;q��u���.��[�P�s��e��L9d�M(A�C3���͛#��iJ��Gأ��3ۇ�Y�Cf%/�+�?ѓ|/���>Ca�>]��M.�A��	Z"�sM|�V�^��"PV�A|-�A`�;M3��O�a�
�6#�;>If�Y�9<��|>��F�P�Y>����@��"��&=�$��+�uP�����'����}�v�ET&��՟�CgX=
S;��,�1�ǩ��γ�1j��ˠL���Dm�Ƈ'�Z@Zf��SI�S�����>���*Y᭞���7Z�W7|d7<VZ��ٍE�[��NŪ����`�pJ}�Z�L�������Y�s?3��Iʽ�
�<)H[����ᅐ�+H��mt �>f~Yt~����(�ۼ{�UJ���k�i�bpi��Mb��?�c��W\ҩ|�z���G"D�q����i�Le��*i�_��
��K���pU�,�=��Ώi=�6�`��(��u1��7��D����9�)N��Ü��&��x^x'��8�6�?ڋ~�t0��q_���s;���Bm\؀}}v�+,�{rSa�?T�I��qJ��d
�i�D\��?
�C}�2��-HQ��1y#�����9ɍ~���A|aR`dx������O�Lm�,�Ae�j���[�ky�h�� n��c�5��&����&~��űd�m����4�ҼG�ڱ�C�ܶiŊP�{e�~�˾<�3_��=�Ö܉a�5MD_���]/�x�1e��B~�ѿ+ح���u�->Z�B��򼌷.���|�ĸ�!#P��&A����5� �ǰM���	�zݰ��� ]���l`�1�X���-�l�A�M�Z���]�5[�,�=H$ǲ�#��8���J?���.	�����o+p�a	X򚭕��q�Lk�y�kY��Ǫ���:ƲE�ƛO�4Ѣ�^W���c���](�ďG�]
w@�C��>Gr��M�KHBCyG��R���`K���,GFMsve�A�ۿTO�V���N�b�q�+����:��F��������PXyskm�^s+��VI��k�$  +��Qm�7���m��
	C�\�l���\��������ŦɨɁ)��MF?i6�nu�8]���1� NM��v����Y�*�Xe=�+����j'$	V�y)1���S@4���0�}�����r�+�*���L4����p��!>#>�O�º%>���q{�M_h(턛�<ި�]�9��z;Q�h �.ێo��`����:)����Oq�-X��²�����?O]�~9�Le�ȳ5Ʃ�}�Y��(��]=�*qn E����Bxg�FP�/�[k����Q��9-r�P�G�l�p:���!n��en�a[<����KF�[J�ٳ22�3,z(Dx���fV�u@E�a���7��7����Q���`�";�|M�N�
��3�AO�	K��}!Z.��S�k��гTx�2!�x�R,HR���?S8��i�r��_�p�GF�l�@���֮֙;A��^%>�%@�/k�T�`��/w�R�NY�&[������Wd�l7�pǾ@��^�\v�R��w3y�J�W'yK�H%2םY��/f��(��E��z�gg���=:��<� _�JOʅ�� �#�ď�)�^~�H�����E��)�PRs�*-0T�@>�AF���*^����"\���u�?0�D"Z��ô_����7O;e��)�d�����ԒSҤ	��
�K-	3�HU>�~ʦ�ğ9�D�k(m�kR2Un1&��M
DЛ��24�b�[Wm_���R<]A*�B̄��T�X�S�MatmL���#<ͬ�`6&�r��C�{HG��%�@�)sF��ʘ�p�u>�Ԯz��Ӛ�1M+����>i�pO�j�=�ў�/�V�_�<N��[�Q��� ��{��BW�G�ώE�{w�lCJ��4�p�=�{�A����A����G���o�JZ|�\4L�$�/���f|��˕�B�X�u��DӔ��O��YR�
�s3�#t*`Q�
p@���ҠfAa���J:�>�UlaNikV��s���V��_�3�$�+�����|�����ݽ5� ͒ǰ�@�W�0�ԙ��z"g{״t69D�\@uS��9�%�5=��j�y�74s�̘Zx�1L�T0�݃�����alqer��4r��"�-��٬΄8>eK�����2>�5?M���mr�N���m �M�|�_��-�!��8��D�s)��Wa��^�d�M��AA��'�5�%��a���^��SZ�`HCŊS����)� ��cpb�=�f~���&Na���<&�)�S%?v�r,'D��iWF��BYgpԫ��(�UoK�s6%�2�w��zO�HFv)����l�ȱR�hT�*��ݡ�g��3t��X�~�%��5��0P�c�Dotg�.	��	E͂!A�Fyfv0��T<-��	"; �?��X�s!����---���X�M��ָ,~���{�0$R��G�+3>V�܇��o%7�x�D!�%�������	�-f$n�̧jz�>]!�.���-�����g_�Gf[?U������%��R��)�0�Z��?�y���ԟ*u�n�Y&qD��қ�o�MD�n��6�.ݮ�LL��%4�Ϲ��Q��5;�Oy���ɸ�?��o	Y��݁�n�B�фR����8���b�8ۏI�q��Ʀ�9+D�3g�����<�d첽��d����� �@4� 9��+���	�!�J�hm�mۡ�� d�t>�Ԑ�1?�H�;*�/y�շ�s��Êc�;��o��J(�.8�*�5m���9��_�j�Ԗ,d� ^��� ����}���Z���8@~�{WqR&���m�Foh̪_�֗O�۫��aJ��~C��d���M�uOĢ���lP9u�N�j�ѓ��&uW}�9@}��� #������øo��I�t��0�ϙ@�:Q��W�]� �g��0��=�,%<ふ
���d�,"���O�R�<B�փ������x��!��EK���i�}���j�w��Q8I���)�^=n��-�.�ǒ�+�I�[;3���bOX�	����F:���)N�+�U����˨ɣ��U�x�+���bj�]$Q+e��K��&E�����"�jcnF*3:���k�I��n"�GV���-~9$-�ؠ�2�Ϻ�]���;zN���x��p(à�� %S2�����B��٦y�if��LS�3��V�b�3�.�nfW�~�Q[)\k��)�>�g@v�&'�^�n�a�x�%��@�/8��dA(j8� PYş�a���/�T΢���Z�n�K؉�y�W'�.�v� �Ğ�S(�ߒ������L�����~����RY���NB$3��+ǌ��eu3��n��O��U��~��i-���&RH`g����F>�x��U{ڲ���C2>>(��T�$`g_8د\����K��l�	���>i����"C_�*ߗ���b��?�\Q�%���d��}�D����h��V�\:j�������\�po��k��p	��BHc��}||j��z�@P5�
>-e��̠7��P�͠i�0�Xj��-�I�X����O1o�O�Ϡx}�_V<�xSMou���`�κ�
ҙ�T���6���	�U�vo�l`�Ƙ'��:�cI k�+rM�b�HU� .�%\,~8剕wu�B)3c {ʕ����7��Z�
Edj�b��<�XF���IZ�m���, e�B,J:4�غ�p���1�H@Nz�D'P�n���������M=/���y�|����%�����@	P~ ��'
ʤY����p��x�V���3�w�1f���g`��Ie6���r����;r^�׋�ʹA�*���!ճ�vy� ��7C�a�Ⱥ����TId�P�Um�$�p�EPt������9*�Lיs?���Ѽ&���}3��(T�Y���j�]��2u��+�Zҗ.}�<����zN�n�^�r�n0��P�'���Ac��� �mu��6L��eF����z��p*� 1i�:�A�endu��by�W��Eg�.���'���+�)�)��W��4]�'����%$��{5�b��ȥ��tD��8ը�I��dt}���EkB�6v��c�y��f]#$̑��'�۲�Qv�+@��0�i"�n�V7��$�RH˭F��Բ��}���.�f*4����P�|�)�2�Ŏ���Z;&�~R��I{��ȭ�~>3��|�l�1��o���C		s�<z_̮�kI�t�:h��Z�އ�ox$��h�{_�3�����)TNY=�/{��e�49���F /qk�>���kD��I���/��h��������!ڒ(���Dj؉�R�cr((���+FrkSQ�s3vA(4_�����r?f�����E`�U�vh)A��"u�-�^_%^S,���l+�#S�s���E0&ޓr��ǌeQ-�5��aS�u�uX[����g��ʜ�1 v�e�����`H��F�����ꇌs��猔+���4�X���F NF`e�
�W&�,@�P����[�>CwMw?o���Q��p��Q�%)���>g�^�?���1k�m���;UWY��US����&�2:���E�/Z �$�9$�1Q~�2��5�_�*�)}���<���y��_��u?l�M�cu��!���$���u�k=Ǫ�c3���,;>���0 ٣/�T��[1� ��ɬ���S9ۏ�UO�~=L_�r��: q�l�����^7b��k!�m��!��C��z@��h�m̕X����|�a���1��u%tw�p��U���F�9l0]�@�-�~���<g����G�K���<���'zz�B�e�"��w�J�d�B5{�����}�m�V��;�V�猎�8���~��Qɻ�� �#�ުΟ��2�2���!�5�ö��TA���p��Z�j�%���-�z�exu��q��,m���t$w����%W��6u���&��ă؉L�zd烪�ϱԅzf���nſ�G�揵!�:�u.<ЯϗH�~�sX O���~ɶ��ܼQZ2}��U[�B	4�&�<{W����D�5"$��|=���`�O��d��Vۃ�ڟ�w����������g�3����bnׯI�٣��:T�͌���I��M�5��D���	��pը�. �a��Yo�����L(j�M@��]٠:�o���Be���2��9VgE/2��i��)�3'��2����������жH��!b�uݝP��v�V�1����Y�
8L)�p�����C���  �:u/�+x�s�:����b̿3i8�>)�J���}��G�7?�g�՝L�_!�tN�K�ʍǜ
�|�>I�:���r]`��;��Ҵ��S+F���b)�	�"��q��_6/�����R�3$���MQ=�7FB.'�������U
L�s�\�q��!zФ2j�d�-k���G�GB��GF�k}er*����'-�/���F���ն~/j��587s���D�l��	�����w����9B�����I
PJ*w��?�g��*2%5��|K �k�~��2̔ҬPS�M=ژ)�?��Yiؠ9���$����i�a������]����*U���c	���`�EE������cWْ9�,ଓk���gq��*
��b�/�Yކ=��<��s��9�;�	�U�/��]���7��K�ȟ��4����-�aΙ���TI�ge�̛�7���,0WZ��.T�̴����Ta��	�Qvz�+q���A_�{�b�����{Wo�t�.�4_b�}|��IKƕx�1� ($��\̕�
����0�!շ��d���m6w������1�j�:X�J�������5��Qo�K�l&�1U��/���`����Q�!�����o���Q۬�䚿T.������YHs��6�,�f�kiZ|��@���9�a'q�?�����DY�ʧ':tՍZ̿R6��ۛ��o�~�Y�sb�E/��VC�6�a�fv�G��myoW5:���� q@�,�cL���4��C���(��N?\<�L��p����/������$�W�;�n/��ɻ�^�[\5,�TX�'���r������[-/��rC|z]�M<���cqp �DU�[���m�"�&,z��rH����<6��!"���c�����|�r:x�R��,0�Y�y��k2B'�OgQv%��5u���.��by �88�t��kA���~�\���>5��*ޅ�eub<3��*7@���&}�g��e!.�a��-�nت $������H۔�T&�x�۰VV��2�Uy���ͫ�ХP�q���<'^u��+I,�ەYV�ܭ=��KC x*R�=���=\ ���
CM
�ņ�f���+a�I���gL���=S�tj�w%S�0�fH�X+�;s==?��o�"��
W���6::����ͬh�����w���Ӂ�hO���&��}S�~���H�i ��`ukU�DA��5���^5E�t�@b���I}>M�cɗ��6;I��kJ9��E���6&�m+��[��)�4^!7�T%U���.W"1�B��zQq��U���96]J�����z��e��R����]vԜ�/� �,�0����uk��f�L,�v�:�Lp�E�0��rc�j�~����g ��� �o4��������x��E�s�fR���(�d�j�p�;��m+=%zBܻy����a{�ӎ5�o���9��@Xun�U�T&f���OH��ćH�n�9��������)ϕ�6c�Pҫ����mW�����<<`<����}FN4����f�Bݘ�?��Ig}�*�@V�]{�S�N�<p�n�`��p�5D����|Vq�U!���T޷��g��X��N�@����@���g��BA�\��-�֤{|Ħ�R,R<ejG�kM_dS$��m����K�C@��<�4��ʎ��י�[ߐ��`���7ю��I���Ȃ�jwba��L�����B��w�(��og7�Ir!����M�_6V�gU�"^�@9���1��sq VZľ��$��H�g��a��`+ ��=���o����D2r@f*���}���^����VYez�_ө��w�(8{)kD�v�)j��Ձx������X������m�j�3G�����ETuʼ��C,D]�>t;[b/���•)T>�����f�:�.j� �Ba?3���z�v��Y+�.{�s�I���9�U���X�V�������f�2扱Q� Wn�	�����	���8w/͵Z�p�� -��X�˖��;�Tv�*nI�#�}�4��d.	�O_�f�.��3gd�,SrU��`���U��f�߆�*��|@Y�_���Q�.�ncw���P"�R��I���9"�֏�j�f_�W�}����"�G�$�ťu��&U��C�4��KI#us������������?��2�[�a 7H�\(�/�#G���3�=��?���b�@A���������t�*6��B�wfHH��O��m{A���+(mj��o���^�e���8.ƫ�bu.a�D`u�J�o�I��u����cRm�G���[I8Y[M�$�m A@1X�/t� ���
�jr�@f�s�溙�6�t�«�7O�Գ5!;�X,����ѣG
��@�Y����tC{�k�싞9.��R�;���ZheW��ު ����� �}S���Ɗ����&��-����I����$7�����#<|�;��ylϢl�A��˨�P�wݲ �0��ƨ�7�3�+�O�}i͸+Z��k�aS�#�1?��C:p#�;s.[�~��{[��U�
Z��_��C:��T�R;����P�7�X�
���q@�T�4]<ؙ�0��v���|B@e�������C^�5@w3+�'����10�����d{#iM��a��
���2� 1B$P���NM]��.���7�� �634ut���L�,�v�רoX��g֤|'n���[���̛����1��?�>&�|�=D���ҝ�6��GR�Yb��0ӇVQ��؀w6�C���ʍ�x�3�-�BBxvTSě{�``��vkp�Nw@,��)[߅*��9K� j2:���Qr�|�?�O�P���r�.A@)DOz�Ig
����"t_���u�Y����X3��*��h��,�������!��mF��.ޠ��vz�Yp/�a��J�a��y������Q��U� �#�>�j{\���|�k��`��V����V΋F,��%�s迖7�.%�����PCTn����QrC���FTsTZ�ώ���� �� �i����yglШJ�htN� �-@3ݒ�ְ"��8�o����@6��r��q�D�=�"tHIKd�xC+?�EH�N}�z�a��"����)$7Li�E�� �P+jm��,au^��w]�x�f�C�����ߗiD�BV�H(t�����]П^R�)8����ʢ�T��)�s��(����E���.u�]qF�-I�Ӥ�OԬ̯7�L�Od5�;\!9NA�ꃱ�9�'rVhe�>曯Y�d�L�Г60$���5��"(�����j�1T������d��FD�Aw��z�=��A�͢1s|��w�W�q���kc�G���^��}�����AWܘ`o�p���Y"�����8%�7[�B��������i�ùc?�a�ԁA�vF������X�qA�G\�+�G��U2~T��x�(�1�Ϧ��ag;��f�sEZJ����]⻥�h`UB���<�'��M_���ɠ�m�JB������v��L"g^��k_g��-&�9U���`P�ZBj���}S:�bG���9���B2"7Zf�0�0��۸W�ﵽ@y���6�e����UE.8|j��1�ā��x�u�=,���V�8����aɤi%�q�8'x��",�s+���6���O�	�\��)�$� �����wZ���)
�xo
���I�Cpu���nTܹ��Z����׹#2Ū�]1ߝ�C:Yͫ�%��W�z�J�������$�B��x) Ί�|A�@��Y���i�r=VE�x}�݈MD�������s�$3}��T�
%��f:#�j`�E�A����>���	�����ٚvN�O!��<�#
�g/����z���y�ޖ'C�U����d:jlDʊ3{ǭ��TAH6��� �,�rX��7���#EBh���
�gDU3���w�T6��I*X����I�Ë�\�s�,��[�� �!�.?h���;)�D���u�m\�H�o����ga�?��-������J:�����'�n׃uu���L�RtRy�2/�<�>p��!���~�|��݁e�Ȼ��e�������x�CG����M�#��^=o���LF1��X.i�,�~�
��4�x�	؃R�iq���z��;G�� ��u���i	���������>S=��(+�J�=��i��뉑~Ya��D�½�rT{�0�}�~~m(�7�Pt�_R�c���*��K�FR1P?�
��z�G�k��6��n�V��9aP�"@0�&��f���w�|N�%f<��+J��� H5��~��Wg�q���Pb����/����ٟ�S�ed�\Lr�y���>��$P�ɶX��r*�a�o6w��-����څ	��/�k��:���Z��awЅ2�2�B��@�4\�o':�QO���Np����R7C�����{R��;�6���s�\�/>b �kË�ىb���ԨS�ж�LZ���X��0��hQ-�/�`<%�_�D1�!Ѯ\�;���KgE�"G�,��ƽ��p3�~E��m�p�(�ϩFF��P�Ø�qB=I��cz6�[u/�Ս��0���\�5%B ��_*�T�1WK]i��G�%m읈�:~��U�wk�����>�Z��Nb(8I e~0뽢�<�r��N�;��{�a�t&hI�b�+%��S�"�a͏�P��]�t¡t�P�����`k;��J�.]��`�ƕ�P�h�GF���s�)r��K�2�3{��i���3�D�9ɻ�%�_����/��FŴ�u���T�ZW���Y�l1�7�Q7@.ôsU�hk��G+D���>CDD~B#6�� ��!Y^AB��;����Υ�'�Kն33�����ѝ J 10�#�&'�g��VXorcHR�	���p��(6+���V&����+�5����gR\��Յ q�v�u�"_��p�]���)]�������s�`�[�0Ci�������:Y*������P��l����&�ͪ?�0(��K�8{����FڌGc��S���J���n$���O��ߡ,��}b%=�u^����#gB�8�2Z������(��v� ��x��I���ڐ:�W�|�}E3�R�-����s�����؂R�W��L���Q-Vyٯ8洘�F��l�[Zm�r}�͍^�]����a|nPcy:���նl�Q��f{y:v6�n������J7B�������/R�ݞ+�ڋT�-��;u���05m�	��t����j
G�8��F4�5�˨��M(嫆t���9�X��ʛ�a�K�ҍ�˷��A���F��ETG�Y�'���ll����  dwv���`p"�}���@�X굝�^� ����d���ɛ��+8\q|ܡb�)sW��7����^�&�Tm�v���h
V�M����1�f@���]�����cB
H>ϒ3*����
��h�^���-Ê��OH�����j��2Ϗ|���@{�Ct"��]� .��ᨏ�~o��y����7��"����1���Rv���]��MҀC�.Q�Lq�>b�o�[\�?2��]�+�I��髂�ͽ�:��|��Ef���ځh��C������ה�8sF�@�;����J���/5�L��%l<�p�t�Д�G�A�y��H3l@��ۛ�
�c1�>���t<�lq̴��V1_� |6*��T\��0��}ƙ0D57�[rj^b]�Ps~��<���F��n(m~����Լ���10z��N����gpcBfT��j����_��T8�2�<���%��	���K>d�I
0h��?���ä��MۈUf������yB0I��*
H̊�K����K��E?>�h36�FF�}�,'�A���wsrE�B=�+�!���Jd�\e(�h�TI�}�'���3O���/u��b?s3i�:U�7~u��e
_��˒�b�{�1���q<蝜��h�6I��W������R�ίzb�3bŅD��j�cy�`D#o���P����s�iE�%�����Y����F6��SA)dC�c&X�~�D�1/�������]�"��Q1_��i�l�
�D㤘[��UV��g`�~�������R�v�_�=˜ݏ?u4O�4S^�[��uX!L�V���ݨ\�m�`GyRwn��!'.ﭷ*�z���a�
���8�`lG[�5�*t�:�y��G�)�>�v�<Y�Y~�	B���Z̖܃[�C��'��&7iZ�c1�$P��(F�ͺ�YV*��QWV
��a�GE.jL��XCr7����S�������mᥥ���9+;B�F5����(�@�A��F���!�T6`4g�A��iNp�������?��3v�����ߟ���xt{��D�=4pr���r[ɹ�����"o��H�)y[~5�9,��f�T�A��J��9�;Si�I��7z�Gh���s'!d"��G_�P|��{[�fO���Q z����Vp�������YW��c���X������I{��=D�d{�~7W�^��S/���	{,��Q灁iX�,X��u�9^�|��e�{3�}k�2��e����@�im�^f�y�\�)Q��c��
�Z�s�J�n�x�.�2����f�?�����Ј�W�S��%��HM�=�ܹ.��������Z���>�B�UK��=@�-��C�0���h�H*2d"wW��q���'�^��Aa���,�(T�Zn�>!$w�[�2���{�����|,h��or��\i�I޸H�k�'�4���؅�p� �#|�r���j����|��9x���~������h�A2�XT�T���uO�mO����� 6��x�z�)i}Q�,YNUꙂ	,��p�����D��4p[���#�R����
�\p�;D�`��y�(ksOG�ؐ3i�b�=u�cց�g��v^����ʚ��Ow_��U��E��AK�|>X:v�uۓ���],���r \����퍯�<���e�u�q�9���I���5J�J�(��V~_��6�z�޸�e9VoG��l�27x{��!��gh����"�]2�E�G]N�T�dK&�M$`UF���`���u^գF.�7��O����wj�z��u��K����frB�.�]��������,��f��x?����U	���M�#lmT�oM��$,6	����у��3�4	�;�(Z���^�Z
����� ���[+�����+�Ëd*�m#P	�3|'�v��힟HR= 
+J&-6�
s/x&N67�t@��i[)Ba�'�{`�&���qo�Ҕ��;����O��07�v�.yE�{��W&���-��t3am�h� �h��9�k0Irr54�wD��Ś���*4X_~��ﲉ�BI[lT��4آy
��PtL�dh�pK0)զ�0����ɏ!u'�$>5�D-s�@�=ՠ�#k4�^d�F�{��F��m���,hw捌�Ri��}�N�����s���]�e��Z�c�mX���Uf��\"P�O]򠪄� ��xӶO��@K��EP�8��O-��.�7��[��b��s�m�L�_�B����B{�3�w5��W"�'�"P��1�]�a�&��qz%�Mc��F��۹ϩ�%�}���`!�g)�[��CT6�|a(�c���&;�fzB����X90z����4p�j���B��a5ἧ.G�i}�(�F��=���E�HI�{��Wߌ�B� �Q��(?�XB�� ��WT�$��Tff,��V��@"ܟn|��f�껂f����SN҉d5T�0�	�شG��Ki$.v���g�W(I9����q���(h�����W,*��PR�|i�#�@���J��ܒnk�(Ӕ �z�'��ZM�w~PDְT�[�?b �5���<c��}F������y�?�8Qn_�;�i���'_RB^�w���{� Ũ�C<�6�f��kdLz�4xG3Y+3�\0 S�FRB0��P�=P��a"��b������u ����X���>�	�OX��(2@١c�HG�D�N���fU4�b����$�:�t �p�oM�У��摝O��7���0,�U�C�kӵ,# B[yNi-��4�A�����Gw(���-ΘzånoCm�c�j�%�"q���h[�;S���lL��9��� Ɋ"V� 	 z.z�
#8��3���%_�b���f��g��8x��60nŲ�	�v��r�z��布�3�������YO`V���c�x�Gjx?��^���;��Q٨�z�x	�?��Ѱ$�Ω��L&M������)(����F�~��:��jx�d����cA}vu�5�TV��50ɄK���R���k��w+*����M[}]�W��ۘ!�)Z�W	���ɽNԐt�-��������7*L�LaA׽���m��k,�L�{b����dl�p��\?��]��.;�L	a-+�ed���ף9z2M/������1���X�ؼ�҉B��X�@�������o����y�n/�އ�����T[��t����z�����L��S6I�8H#�G$r�j0ٵ�k�p�G��4y3��i���9_���]�7
VѤ��o�k��K�
~�*C�Uy�Ӿ�7�b�\Cb'fi�0hKWB�j�z�!��@q3���#);
�b`P��{�}��QWo_�x(��*||;�S �h��S���Ck����k���<����a���!ږ��kSm��{�]�9i��.0�D�����sM�	P���E�Mzސ��Wz���Q5��ż�Bt;�
Q�4:����]��6LH�FTfO"z�� @�m��l�,]+2����;Nǣ1����B��{T�9�PsV� o��7_9��}-��T��I��:a�6�=A�.qe~o�h9NX������wL�2��Ӌvk�f̬����b��B�Tݕ�;��Za�%�p�!4^KK"sw�e�@��#{J�o��6�^ΰؤ�PDί��"ŷ�G�����J&�P�G7�%��M�i+6�u&=�pi�W4)O�nZS���Z��(('$�GS3O�pn��`+
x7o���U��4����؍K{53K">偵#���Ul����8�0���b���>�������Ͳ�����{cݮPƿ��������⶝~���NڇE����Tv��(����N���}=\B�+�i:�k$�z���A���Tw�Tf�K�� �(�-�:�|��j�o�����-2�	[Xߊz2��c��s��(!(��%�̃:�ɓM'k��N�w�� ,��4*y���9�tHpڒ�Kh��P,P�j�;�~�z8������}�zf�z�P�,+HȂz�p��:��g�	Zt�9?^Gi�f��/;�1���+F���uAq���iQ֝�h�ͨ0��*����c�t�la�?�BH�J��lb�u;ny�BT2�ϛ0�T΢�J�F�U2aK۬�� ���&2&���SC,��C��eYp!��C����jZ�"ݿ�3��Ù�1x0B�ޚw� ��M��Ð��)Q#*�%M�f�˥�N�ڎ(_xaS����dȎV`_�a!���pf#k����xm��Գ_�џLl^���M�vuJ��v�{3�CH�M-��&�9	
��ͭ�Ȏ���G���z��#��V���oY8��L�VCl�!3� �m�G����7Z��Lw�m�w&�6N���Qh�V2sD����IdȬ��[q�ܞ��Nm��6逡��4�P���ܺL;{�R��T��H���nu�(ף�U������i��yg�f����'M�zjX+�Qj�:����P���v��"�{�sIߵn� �$%D�%�N�kBߠ7�>8�mo�P!n�DНhF1��Sҭ8��(��R`�O�L��bÂ+ԕ�a5�$�\�Nv�/<�zM_If{�{?�@5ǋ�(ӥŊm�-�}u�C��z�缤 ��G����^	�Lϲ^�8�{l���oré��2��L�³�rZH�`�%l�����t�$x��C�%�?��*XHS��a�b�'XG�£�U�����Q5���$���߰U���̏�-A���V-$*vϕ%ss���p�D��������cO<�W<
"NE�h�H���JL���O�ݠ�	8��;)�-��4�ó�a�Aˊ����$<E;b��^�fp���9;,���r����^�'��8��O�(fwI���y^�CKhHb#:o4VW(J�+Z�NS�)��r&3^�c�4��+i�Rb��/�õ�� jCp�-��?�#��;U�'~� Z��~T�=
Hڞ�d�I�!����.�R����i[��)�>Qa�w|���u���oP�K�q�ny�^:��ׄ3��$�HL$��9��R�3ə�AT�,�?J�\t)�E��2Ӆ-��i�GS�#���T ��!��x8ⵜL�.�&:�*��x��m=t?�W�DK1���I�tP�1��t5)$���Tف�Y��$���c�M9� 1c�;q��Į��o�|Ԛ�IhN��Y�	_R�vUT7|ͮ�AAS��Y� k���ؗ0����:�_�U4_
��t~�EZpv���#��?��,��M���*��j=�~0?�`���\�� �,��[���{B`6^v���l�(x�I>���V;^�S){�f�$���{ϻ戮�~ᶓ#z��a��綐~�46ob4+���X}�>�`G���Xy�`�)�,5��������${c�{9������y������Z�
�)͎��D�1<Q���@�=�g���r:�m��%�p��$�y�R��Q��B���=�"����ҏ�2M�����+�#��0�w��ޅ6|C�f�lx���������m��p܉�*�f��&)ʸv%�P>c_taB����z+oI2�B�b �a�
#W�݄�9�g�Hyÿ�%K{�zӹ�}y�Y-T[��7��� ����<IQbf�nC������b�=O@�Z%��2<�'þ�j�u�J�s��q�5��d�����mt�O) �:k�{-7 ]{/EC�&�����k�Ϋ��V1�V��8�����7@�=Ҝ�Њ�F��f\���#��u���l�H��I"�o��j��(���;a�&�:}��6-����֠[i��X�/��[�F�����ǰe�0d�]�A�f5P��'j4�8��l�_%����)��؅��hBT��g3���������wq�xȊ���`5n[�/s��n���Eω<���)>��T�y����߉�ok��3i��`�,��6x�܆�:U~
4��tDo%�
�p<�۳�#UR?;h�=M�,��I ���ʧbgE,d�z(9>^�&��;H�9�=G
�7���Mv�}�v��(���c�L�ao�
6�f(ckw?w��QNV����X����o�c�oeM����ͼP��S�KVL�� .8���]�"K9NE݄�`�]F%�4�&&"̈�S��og�&���=�G�)���G��D�|��#�9�t}�%�_K�+�$�Ɓ���T��#�{,�x�~�q�>MP/5�'�4E��ڕ�.���Y�K9���[ ��*]%-��S�,lF���s^��ڃn���&��u���>�\,%h��M��}26>� /��DRqZ���jD%�_��Q�@-̈́(.2�B9��	� t׌ �I��s�&&���/��I`��y�R��U�����`-tӌ�����_�P#�.p�{�ͤn�[��{u2���G��O�
7���)��+�x}�[�r=w���},k�)7��%x��9�2����dx�)��ZP�3ѧ�� �2�U����↋�,Ev}������B�t��9j�{M��1v˱,�l3����8��U��f��Ê��>��0���א�aӄ�� J�!��s|t���Ѡa�DXz����r�܎5��6�4K��]j�+�T_��XP|ѧ	���d��X�b�"&�͂�m܆L�����^�!C�M��:o���Y�9��}¯j���M�v���#K�m�����+}�_���qU�T��F��<Í�}"B�]�-`�q?�BA���d]��WP�Oq��	4�]^�i���w \���]��,����W+�l�v^��e���d}%�O.ۗ���}�[����X)r���J��%���1g�ٴ��8�"nU�O����ӻ��O�)'�����$E]X�=�c��G�jtQ�B����?( }���'}��H�CT�UnWj�����a��1�O$��p�?�3�L�]�{jw�a�� ƾ
�� ���b�������Q�N.���Jܐn�o�hj���h�����5�\h�}�{+-@�"�G��$뗵�Yg9�>@t�i����N'��I��#9���c���C��$�����i��~����*݊��˔|���3N��v�Ӭ��1y#��ʨ���j�@��̇��h�e3};0%�i�APhjf<�27NQ���I@�6Hcͳª���g���"�/��L�҈��L�Mn���o��� �����}Lυ��?
z'�S��L`�/���'����>�����|v�8��!�(�o�c���$���f�/BJ�������;鬜���H,r&�F�VE:�?�E5!�������F`)�_�E��@�"���҈<�4��g]�QYې#��^,Fߏ&��>�K�r/�e��;�"+'���Tq(�������k��K_ګN�J FK4��Bsm��bv�X��s�7#At(
T:*�=����o#�U�'Z�s�=���crU����Dݩ	���@���nT�UԔ�i�we�����"��@��2�*/���'���o8��~��vęT���ڕe�|�{���Ćjq�r�׶ O�#�HC�>,e�57�Z�_a���1�LjG�q�z�C�z�4YP�3>��EI������jB� �l6�z��^�5p3mʇ-�i:��ԅ	�g0�Ge��N���m�1Fs�����]���� �2�X�͝�aG�߈�"L����X�!�?]�^�(��6���vS��gP��3E���Ҥa|��*���Q�����+k�/�`#D�؊^�U�q�����sՇ���?�w5�k��x�Q+�'ql�29ɔ5�1?A�J?�
��*G�Zﰐ���-IB�q��Joy��j_jl�ҭW��\t�iR�Ŀ�^>I��e�� �퉙sh��z�O,tm'���5��&�ǆ�!���]�	t*�6�&3��؝�]�L������5�鄉5ߓ�}i�3ѥw�5���;���>��U]�ҙ���G7}��4/�W|�i��g�>O��:D�v4!�� ��{�}#�)����=�/j�hdB�GK<�
�E�`G�M�-s,R�
V���2��J��<�{�^ŨD��Ł�p邷汲�����
�w4�A7�p��A#ƅ���?��<^�o�f�Fz/��6Z!�%�US�E �L>��qhW�hȠ�)�z��	��ut_ѧ�Ѐb���`��#�/�X�	ť�%{NZ����<,'s0�������)���IdhǚR��M��>t��Le�LpAQ/:����y�i;���`LIaR� =Ǔ��K��Gz7s�'�SWb�4��O�Z�6"�<���{�P�JXB�{:���ŕ��x8��G�\���~��'@����N���R�6FO����BY>���9��LE*���c ZE��7z��w�p$���J���[��� ��6nYa�&#B�V�&��_E!r��4=i\�b,���ɕ;ҽwQr������^/��\nN��M���j���"3�{_kѰ�o�Gf���$�m�Z�Ұ��(�Ϗz�� �:Xb>B��K�uM�c�����<�����#�+�%�!��{o��L
,DfaS��u�ɖc3�pA!�L�]	?̆}u��|b�c��>���ݭ˾d���jψGx���aT�<
|bl��y/��GD�%%�?rŕ�̫"��(t�d�v�$]N��^���do��jܩĳ��ŉu�d�q������Vy�G�}�U��"��E��d^�[�����{X8�;/�]Wy���$�u<��s��jIϻ `S�[0������mOR�~3�"���	��I��9�\(8C�?	��y]�_W�3�x�>%���^Y����쁦�ss��G\�n�}{<�-H���0����I��n�?��m��[Uf���>�[l����}�,�_b0;��=�&�!iFmro����j��7�J�*:z�H��(P�c�:���,́ �	�D*���y��b�:|�Y,v�
��br���E��)���{�]	h�CU��[���Q�T��gG革x5F������z�J�WTˡ����u����'����-�L�Km�fگ��N%��􊃩j���t )3�aY������Mޢ�����۬*Gk�ҋ[+^���'�{��VGɸRgi3�D-6�(�4#N��xP�5�CD�� g���y���.�E众a;sф�^a�ק��o�}�߁�8W���R>���P�K�-����%�����`q�� %�]�4̎�A�&�������d��
�L�N�k}"2	��iB�u���mcF%Cu�b ����O�x���dZR��NUz{��a��z��11��d[���]���it���7�9���2_��z��"M=�%b'o�O�@W�i�����2f5��4ѿ���q:���IW-��T�ݺ�o��6�Q���V+�-{Č��IR��I�Գ|�ޔQ���5��y��WO�|V3�O?'ɺ7_���zQ𣹫Ӭ�׏5�V��"�DW�[��,��z5��y`�d:���Y�^~3�N�]	����Q����4T
�<��E��O\������9�/���b7X�~�����{��������@���B�)ls霸(0i�sg���qTQ���;�U�_�¼�ْhw %y��<׎��>�-���p�A~1Y� �Yw��!�#�Y���>S�^3 �� f-(�J�=�v����#����~�=bl�(��},���n�����
H������B89kΪ�,�� ��;�>5�!b���r]W�:��wije?�p���d��Kj ��o�D�@�k� ��-��`8����^*�7p��'�rm�L�3=
����H��J��=�_
��ÆCȰ����6n����f�34;��ɲ.����"�_x!������p��|kOPt3����냜iN��tT���T|��ڙsg�aZ�][�����'	=F��'&��Jq�x{�� � ���_��$hj��iO/V���t�I��$΀���dX�x�7bn���B�4rx�0�?R��3��9��3s>_{�6�4:�h��Z�V����u�ݺP�P��zEz+��=߇ZS��Z��J�J}��ӡ�ܝ�ί����2�7�P�'�]�|g�8ٰ8�Xح�jo�"����Ϧ�F�)���)���a%vi�����?�h�o~=�����;M�\_�9�̢�#�ͣ�wHY�����Q���8iS�^��i�K7;�;b)�K'�*Ҵ�>@e�#]A~�������`@�q�����l�ڊY��5s�{�s��Oƀ1��!T������W��w	�HA��L���<y�p�!$��T�%@���s��{r�����۷ �}+t�7��#����v{,6^Un�!����j�X�7b�y*��,��T��c���L�	��~�����bplLg�#���A*gtX�&pA~�ޒ��4��e=�����0e�g};5v��� T|�dy2���:�f���#U�;���	�sv2��|Է:�h�@��oں�\�Ksɾ���<Vl���ζ��@��&X���{��̙h�B�B_�s���V���7���@���x/����t"����sb�hկ����?Z��U�q,��<.^6�4��n�h0	�9�����8@�?8��錔�5ҡ)1$T˰&�k�E{��܅fw��=����c
�I��c��3~��vU����(A��?�"j�Q��ڧ5�����Gӣu��K�BB���rDi��ج��=�>��W-�oQ��]-G��5ʤ��L����xĺ�D㹜�T�� GX~{m+�ı_��D���Ҁ{0���f⫝CQx�� �$�ʄV?���'�����{Y/a+��q�wZ.0������q�-G[��7��լ�'ϝ��T��H:��Ǧt�vw�Q���-�W��qw$A�t�mY	,밄���C����c��Z��ܢ���ȹ�9��Qt�R[�@�L�'je逽�OȤ�8�&�(��^Ck
��02,t:�6#El�݌��b�,�����8�ՔM�[�ٜQ'X�z���z�˝!:�k��/[�����XTos+�u	u�3f�V�SׄOBR���\�[�G"Ku\@�p��y\?<�gslQJ���yeAk��$�X�������	Y�7���b�$�%�r
$�m�|���a�:���T����H��V\)֋��=d��XL�ʊ~C���vN��0���&Fhg�$ >�-4��5�`����3U�MEd�ː>�	��U�u�"J�Z2JElk��\��Bwn]�C�^�p��� �9��8aWP9� ����f��|�Tp��8��J��$��%@F3�K��8X��W��˟�[�
c�q�\�z�b�-R{!S����%b%iOϔ�ͫ��˸2d�@��g ���nҝ0$VJ��9y����+�X%W�{�#:Sȇ��eK(0V��!��|~���e4�j]x��u�U&��B
||����wA{�ዮ=��EMx�l�'����M�S�x'G��Z��k��}��Xq�4�=���
>&N c��A~M����E�ax��!���ݽX"��J�8RD��=' ��Nn�9�͂ո<&���"o}B����5\���/��a��>\hV������h@&�c!Vx�������ڪ�k���%�oVw�$���8m֬[ʏb��cF]��;���٫m�7����41Q4��zt�WG��X�4g����r���3*q|Bm[��B��VĽxi7�NU�A�其���$N4߆N7�x�}����m�� ���ۗDs��7�r$Y2�_M|��}�R���JOk{L��d�Z^	Y��ۀ�367�5e:<]S�9ye��bNZ��n6}��oc�ey"�"{�݆���e��#�>H�]-�ȸ�G�Tt�Ş���8Ȳ��.u6�/!��g����J�;[��!��[�m�C?!
�Tcn��S��#]�ù�]*.#��b�������eUc�l),��ˡw㈵�.q�h؝4�3lT/d��;qw"��^���0-�z]��<�ak�_44��]�X#�/�� cnN�Q��x�N��KR�[H�A����cJ<%�!t#�ے.��GJ*��cG�U[�[*�g��N��t�A�^A2]3e-���͘�f�<F����쬸���$�!?/�L�Rz�N�ŪAr��p�r���P���߮��i���+�Qw@JbAЏ�5F@l�R�7$�JV���2Щ�.`}��".�2�cL,|T�� (�]v�����H�ٹr�)s�n�g��Y�y5��6��H'��ܖ����|����5�e�'�`ӄ��*��xwad _%�BQ��Hf����&X�0���|l�+��y���g��h�������|*Wu�̶] �X�ކ�����]����v�Jo�u�]�8?�!�^�w�8a��8i�N������!�O��.��k�#B��@����J�Z�c����i���j)���Zvo����]lh�J�k�⸂ sZ��3�s��;�C�0W�T*�s �\@D�x���:�mh�V�	r�
3���k�p�}u%V�U]{����Ej����(F�H���	�)v�v����&|���mel�0�� ^�.]6J�b�� A�m���40E�W� �Ъ�2h�m���1
��z�7��TA5y/���<t�5ߤ��q�L��%��/��i$%�"��`ȶd�QT�"��?�+���Ōz
�1h��*&p��)���L|����+�h��moʕ$�}�W�nTt����*�![)4)���?(8��U�T�N�,)Q�e�[#�1���2�r԰��I��̈Y��*�S����V���������MgT��c-�|9�
S�\��Ws��~F�^�����D�[` ��K�3l�K��t^�FF�}D��K��yt݁�~���aC��N��q�vr)�t�G�����D{������λw�@���X��g��~���@l���v�q�g;�l��lV ��ܰ-cS��Kx�Z�R��DξJ�"�ϛ.y`�f:�B�����~QP��u]f��+T�
ؗG�bo���I�	k���b�����s����$1�g�����~8�	t
�T=V�qI�,�)e�c{:V������z���es� �X<��%�P�G�ӎg��-6d�>���#P��苳g~�^ɜ�g��z�E����f���ΓU|50}�jv�� ᆗpC�ǫ
�������h�9���G�V0ϯ &>|����DBd}07�+��;_{ �#��Jyv�Ә����)?�)XT�;���?9�~�?}�Ӭ�߼N4���5"dw@~��+�����s�PN�9DdnL�.{�l���7����?e��0Z(q'/%<���T�qœs�E�90��z5��3�Eઑ�t�����ݪ�b���E�� U
��Z�r��2��o�CY�q�%�]��a�� ���3_# b���;t�~6x��/��Jz��)�����E��~�NR�D���a��˴��8j�	��ƶ� ���� $�#�>f����_�+�T�*�����\�M����9�H3���)����x[m�a��XE��k{�j��8����g~�Ӽ�I|L���S�I]��Wq�O�sW�e�������/,����z�D4���s�f7n����̓�e=g����6y-mv�p��mHtn�!߼"�9�|U�f�o�Vr#�����-��=��8
½#spe�I��#sS-��!�Ä,��tl�uҾ�76�O�Q��4�o���~�� �3\`vx�����RO^�m�R�5�Uw��~�~��V/T��U;%O�2�2��˗s[$��hP���[����)��
�c=PJ#�_�(
�C��_h:�
��� | ��=Q���;,9�|D�=D	�������v�s7�5&Ae<�n���o�=ҵ#�3%��Xw?�a%2�/��1!��׍��q����C¬)�ƻ�J�_S����p �܈��V��NyUt?I���E;f�!����� I0#�f+�n�G3{�|9r���ấ�,�R�`ޗ�tp���Ԃ�i�6�
�x��/�C!IE*��5�:C=�*��/$��� �-���%����(gJ�^��i�mC��(J�<���Y|c+����o}E:�qD,7�^Pt�}��eq�0߰���Me��'���Vx:��5�������}~{�Q��矚�����h_�4�N�.�|��e�� Ȇ�6A|b��U޵01Y$e��+jB���y��N��E-����8�嘻g�"0* ��/Ays�Lk��,k����>�n��~?Ck���^���s�����Ǹ�o�����_����sbQB���d�����Gu�JAFg:gq�_	$7i�BP3�QX�4V8��w�oAWʶ���y�VD���;����7���7>rC,|f���������*
)�|%�>��f�l���9����� ��R?�_&��.4r��O�O��>���n�P)b�'���0����G�cnw��Y�?h��L*�=��ur���k�ى@��4V�o4�[�g�X຿� ]��z.���#MO�/���*z����g�#�?#p�=�ʅª����w��r�k��8�/w������Y�ա$x�7�S�f�7B�����6MmgB��-�\2=���(}�2uq�ϕ��0[��tA�4��z�gV���*֗��Pu�k��0cw�EѪ`�F�$jE����"G���ʶk����ݧL�8����^f�3,VY��
N��%�wlJxט�F�wS7Z�@% ��||uDY�=�1�.ˤOG��Qo�i'��d����o��b�n�1.%؋",�9�d��:cK���l�煊V��"��!�����B��oi�k��~8Q.	��L�Z�����Q�T���W]�	�Ϋ��ߢ�GF�\d�_4�K~r�%��FT�Nڍ�	��&��F�n)�u�D}�F�z�W���ٔt*�!`T%����dO.�D�'&�!*Y��հ�<$�~v{��i3_'Ӟ�E�y����:>KT�wY�G	�o�����VW��b
XXz���� >2ױ�:��� 1���cfE#�{L�g��/8r9��% C���ߎ��/qF�F����A�.�+Y��T}櫼�Em�
O�G.��hq_�W�\HA�P�(������+@������Ƴ-{�� ��6�9�:7-�%{��9f���v���h�qG�zE�:=�	�8R�nHQ�ˋ��S5�p{���l&�>����~��ܷ����0H;�g��� {��2���ri'.g�sZxo �+k�ցv��,��wW6�o��&2�*W����u��Vژ�KM1F�兝48꟒o����
mQ���OHN�lޤ~�ʏ8C�!�������\�duɈ���=q5���g�=O<���r=<Դ5�����_�o��k��YR�|�ç�L;Z��^�G��;�u/�J�{��	�D��w�w	��ǢS��l�,����vr-av^	gX�,�5�B�n(~/j�P�A�N�=��i��4����	��U��E���3F���w����#�Rrk{�r4F4���j�\itTiv�?��Q��d5���`�L8~D�� ��������G����5�^�Kq_�
�hOxنs��TGY�=w%5eĶ�M
����v.�OZv�@��>�
��nֲ�t�q�R:��ں~H��t���ᨤ�Е����'��0��в�S(��(��ϫW�4���D�,����g����׍�0��KŘragu���{����P������ ��0��p|�rYx����������p����w��]�2]��W���@�A�#��hъ�Rq*�Ӱ��&�B�/�CE�c��p�狳tG�Jr���U�']G)��`/Չ��sڢA�6
z���8��Om]�j-qh}'=;�k�.�c���Q�.��.�kt���oq^*ۦE(�����R��(t�g.��A/X�,��M`A���z����G�DT�w+q��X�[z|�K��Ѝ�I��H��ݸxH�h�5-���-�>`�L�7�$�5/'���o�v�����^�:���*N5�;e�z�b��^�-����9�,3�t��w�^[fI����A����P������D��&��x�\��S�nWZ{�α��(tl;��V>��`O��J������>��j�z�aeM��G���VZpr�PQ��.>wN�@Q���?��)��@��:�:���qV�n�Y+�%1 �����f���#���%�j�V%�@���&�TgB��]�B��$ݧA�a�N���.�w��Щ1mP�Uz(����Odu���6R�n�ĸW��ê
u	'��a�l���ͦ��{hA�HL�����}]T�φ�X�غ3%w�������`��	ek�S>�5����wѩ
y�6w�)�Q4�I��Y�RR2^w���V~����R��7:-ux+��x��Bb/R�X�^�Οm��[>��ߜ��#;������/�ڞ^^�{	�䭻�(\J����f�0o��T�mZ��R�LmU�7��~:{i��_�	�ފ�ro���:��k�$J�8��SA����,9iV|2X�. �4��T�Q���i�~Lc��g[�x�&>Z��Le �5H#���?ǈh�Dy�.(p����^#Z�{��o�SFC����v��-%��80*9�ڪ|f8� t��+���G���+1%�ǅ���ޝ�=,���:g@���A�Ŏ1�kE?�@���U@'��J�b�� �`g�9Z�|���3hҖ�D!�>O07��"X9FޖǄ)���2��t�"�^�h0�J��Gc@PSp��vۭ�9��]aK϶�p�'׭㬜<=���ed��K1*b��O�rn3T,�q���2:��yq�\�5`R�9��i]��#}�m�;��6=��~0)�r�����:�AiX%  �� �5^�0�w��5l<L{��q��C�j+�$&�dd4�h;�M&�""uL��Оƨ�p�U��*a��$��ߴ�^K��L���($PZ����\�,,�n˛�t�1<�p�4f�>��NR��yF/wS(<���eS+��D��?�r����&N}�UF�0��o��f��J��I]#)S�����k<�P���z;�M�������8l������3�wnX�jiS��Vt4�,;����6���YM��I{Ɖ���f#���o*
�e������"U��5�U�v-�?��Xgg�8rMʊ`o�m���&a��N��4��34��f[�ʰ����l[��h��:���d�6��C�i~�M��f�i6�6�WWzq#{�� ��e�=��T^[Y�ɞ�����ݢF��]���^�T�bH�F�.f</�FpQ��~D%�>�a�1�G+��{��?���ru��%΀�	t�v����;}@v-�f]Sd)���I*3�Et	2F�76L���=)��#����l��w�6/��9�Ի�öK�1ﭶAD�&Dx��%�ѯi%�:2-�[��;��s�W�"?��{��g��]��6jmϥb���:��MmZ�'!gg#����}����"dIOW��?>�O����I�B�0k��\/![N�S�S�e�w,l�x�D� 0D��K���Q�Ӊ���E�M�(��.����w0�m�.�\>����T������ₜ̲�.�Ý�o�n9����0>p/�v�����E\|X�.�ErK����i���-�[�.3���E5�<@�t��2��B�_�_���}y_���XTC����C3_��c�L�\�����L�G������]�`���^m@Q�V��g�7G��[�]DX=�q^t��r��5�p;�y�y �D�m���q	��+�!]����2�ge��Ya�@�s�x�Xʕ���3�����|�
`�Z�oB��PuC�]� �r@h�Xvwr�4�B�;,��s�b��7�#�������{�)�<�%������f�݆#�:�n!)e�e�����_�O�*SC#nSO�w�A���a��;sj�HjSȿD�ȶF�ײ�n.u��������܇>�`�JJ>'_�)���ִl�D���M�/�"3�1���Vu�Ϊݽ�ŢNW�A��
}x����M-W��iU��� ϔ�|d��/n�mz̽_}�qmv������)����ūp�N�?�K�J�
T�)7��܍��x3�p�f_a���8���lqLXoCә���l�]O�_��څ����U��UY��	H�ѽR�@A�Ię�bT_�s@�A�A�:����Q��,�J��wxu�tw���e4r�*�-��X�'��B���Ixx�A���ɴ��H�0пF������/L��譸���0�=�X�3g��3��E��5r�
�����k9B/.H^��X�۶���l���G��p��l��sm�����$�A1ibrz�)-�Z�ƚ�f�r��{�;���do�/Z@�ldDx�"Z�(!n'��,��6�P�,����{3���� t�8NƸ2�<g�@��4{����i. �ZJ]���s��,��E�S�u�T�9̂D�U��E����8�(B��JY ���!�u��zk~�8h/;s����>��p���V{��m��n7E��qd���o�Y��Q�/l�K�8����c�\�h,Ǚ/�B��:��>Xq�[`�2.(L�OT�M��xk*��rI�
{��8�+��]���j;���#J N�����؀\��<��:���ąms�Bp����m�to�y����Ǚ�e�܊;��d�uk����!�9�E���A�iގ,@/����ٟөy�u݃�B����9W%�ķĽ�s�h���q3nܩl 3�-dTpD��]��8��}�tG˵�57���U+I�ͨ:�MĦ�v1Ub7���>�� �
��ԺӒb�_Qm/^+�/׆&�;�#&��TyL\�1̀bh� �'e���kEQ�j�P���$����߃m>���6� �cM��[��#��s�Sg��"/�e[��L��v�_��O��Pg;˲O���| ��y�J�aH���?���%DJ��(���A���ì����dW��wY|e��o��jB��s�K�-l�}�[$}р�P3F����ݮ+��T��j�$�,�L�?�6^X�mNZ��C�Ě7,ht�3��@�f`�h���md�5~v��35v�<�y(�(+,Xc/\�U��+���	jhl ��:ӭ��0�ъ�P��30�?k��ݞ�0� �}��l��D���4�e�����^q��YU���
r�<#ӛO}0é\[+��P��E0�7Լ���q��Aj^g�1E	`��VQ)=Ym>���X
�أA<�dJS��+��D���m�%K�m���͚�tN* �c7b\��mRw{�q�ǻ��U�R��LB�&�'��:�X����%��� ���*ؤl��
�?E����SP�%�A���G"�UJO�σ`),�U8"3�����9�x�
��'ZVb&��j�Q>O��e�Ⱦ��O�5h��s�w������`i���]�[��Pit_�ʖ ���̵nA?��Tw� �]`�J��k�Z���=�F�^�D�QJB�: �84��|�r�>�q��ȥ����O�'tT0�������!�M.��͈BC���"9�5�)�Iumk���	q.{P���`B��d�ZmU9���>O',�\����"w��i�ͅB����>��θ�uQ�U������E:D��ԑ�Wֱ��Os'e$��M7'�'RB�o�o7J��c�_;�U,�Q.D��ܨ�\`(�LF�W���t^��8�s�����B�<J�8��zeHa� W�ݎv�_�g���������h|�[���/.>�·3�
h%�]Z�G/|���k�Ƕ�e�A<j)E=���d�G�6�9�V_� mB�9e7�zTۨ�F|���%���O��u��M�Q�8�㟻���:G�5Wr"ڧ��T{��Y0����v���[�SF��:̛�9�	ǀ�� {�!�cR��G�nѿ)c-�����?���ss-w �@VNR���k��S���Q��&�]G)��N!>�#��<��缎W��6��s� >�k2$��$�f5fx�� [�ޣ�3�t��0_��]���a��ޟ}S�+ؕ�?d�g��s��4Zɇ}Ȳ�V��+{��+
��%����]��9����,s�`��8�U���'{��ŋg���Fَ�:��c���o����o��x���U8l5";
Q�Z>r�����Ԍ�烆&�O��gx!?���aR��˟9���RG��q!������p�RV�6M�^��]�e�]�{K�'�PB���!��Wp��i4t�}�a�g�Ѕ����8?�U�R�$z�D��3���QHz�p{���~�F{ˡ�c�Z�*4֤�~�21�{�M�j��`���P��Yl�T3�������ڟ��a�P��Do�iF�{J���47�lm0��$x�d�Q�+�^��[``�E���f�������"���o�ե�Y�G2�>D_ �+�{i�W��L�m��f��t?���=�$��`��z`���`h_����> ���e�`.��-������AW�S����:��2[=���`�rTj�����PR ���\���[�y��R�k�h���a6����4\;�JY����.Ȯm:5 �KŻ�	�1$��"[Zh�ԅV�޶�NƖ>OM���X}&F����+|G���,YT�~1k�$j�_����M���= �B���ēV�L����j�QF7%Qb=</3��Ʊ"��|��aA�����r��^8[:f\�����h��!כ^�_��p�zC;��V�k#��#U+��7p�\�,���%`iކ�Z?�m��Ǔ�Z���W�x���HwQ<�����k]diZpO���/:���W��ݥ���GL�3?渍�]0f�)Q�n���D�8ZI��q8̏e���5�R6��j3���S�$Y��!3n|B���Iqo����[����"��Ξu��o]���Oj�0�h {|Y��w�&ګ�x�qo�#�v��u������ ����7�dW8tR�0s(��Q���=�~��q�1��#Ɔ����9ca���H�D����򎜼H��a;�O�aOgKfb���� uC�4oMo6�p53<������T�'����\K�O���u��O�\��Z#l����@<ƾ�%�Hx�ν:�b\,�PՍ����D��I��=*�)���nRʶ��*����LHCeǪ"=Y�y������LRj�1s���'�z���C�N���}1����Nk6����r��m j\���"L]<���������-'��tJ�6l?�^�m#~h���i�*��a�L�L� ߉��ÿ��r��0>g��b}g�ԡ�0��0��`����{�We6WI>�_mO�S�{U����m�/|�dC�>�Y�[��Vݵ�2��AZ:I+F�@��9
!��[�	ި��?�dNy��p��?.���@��5q4����O	.��e�ʃ�^GA_~U��xhr(Y��У�d-�q<;?��,ևIx;�A����u����?�����D��\w�+*=­ucty�M�hfo*`��Z#���/�n��Ͼ[,
��ȢOkX{���A��~[&���ь�"��{ϔ�;[xъnX9�]W���=�W|�,��tm�R��DoQl;������td_�R�쯓+9���	+�:��R4���03rV�EM{�i�r���]�����X�zZ����	�U��(�g���s+U�w,%��jj�
�^��I���+j��o�N��~-I��/���fA����/��v�Ǡ�	��I4I1�̠�b��	W�?� �`��������Lx*;�l�ݴ���<������W��7��OK���}&��T.?X'̣�K�~��:ȍx���@��v�n5��ܘ���_8:���؁���EP��ܖ遜��q��ZE� 0��\��N��$��i�!���ȼyAN�#'��D��`5[���S���M΅b�C9_���o��|���K��t�.Wb�^���ୱ|��Zmχ~�d�����,(M1=|��1��ѼR{c���|��F�-�R�#���o����{�����m���Q�c'��G�0�z"_�F6��nf�q?�{����Xoa뇿ۺ\L�j��1y9�ɧ �����Gx�55��6t%���M/�\���l��"�Wt�ps_xG|.��2ӊG-"�f�8
�V�Z�[~=�Q.h�W���3\z�%�Z��%�/�G����㩣�%}��O)�&�0X,������#�S�^����R���=c��T��Z���ǣ��*p�tw-N����]d5�W�#������?�0�V6g=<%�O��a##.�Y}�wTtΊ���zm���]�lLh�*Q�EG�A��O�UWf�O.�˷��(M�w��_�R
�����	�k������F��^M�s&!��>Q�tf��9Nyw�&3K�� :�p�2t�m�r�q%���)Xի��u�N���#/s���'�T���l,�;��ǀ��Ƴ��8����	pII=��T���s	@���Se*�y=>�S��W�qs��Q�@�Ѩ��]�tG�
����
�����
]��m|D�ދ��H��yڑ���8L��:�^	j$5�Xg�=a1 �����F(+�}�ǎ�lRʳ$��\�"��J�I�|��=��sk��c9E��o���$z��Ș�e�E��͑�HV8	p��E����v�pJ��z�ƤjS"aNh�pD�e�*�жJ����[��^�h�@�Z��{�ZAզ���gu����m��6dŜc X�5ً�fbU��
���&O��Ӊ�n)�3�0�C ���EH B�)|K2i����W�d���A��2���k����B��Ǵ,���5�'����Zp(�jR�c���am��o����O��k���3f������)���sv���"s#<�Ƥ�����5y�2�NuW��g�`�'z�7��۸cמ��ߘ���u������]� P��;���4ׅ�u�0|3��ǩ��$��qH9����`@��L�#�j|�d�Y��kV��2����à��=0��ܲ}j�ꎈf�-�>ݝa6=	�b��AH@5���:���soӥ߫�1�(�� 쑨|�k�K�þb� Rn���TM+�Gl6֕�+�|R1�=�&t
���*܍]����,>7�'�F��2SML�A��I�\^ǌ�d�
�J%~PT�{��4;
��ǃe�3���*˂ׁ"�3} ����(K`0���g���T6}������+It�@Dt��n/>e�SC đC�e�a�S*i�-n�+@=�U ��!vs�OE����1�ĺ�e��毼��˫��2�Y\|�����W����������`�d��6>���?t��Fj��Z�ı$Тw-����.{?p-̗�w�kc��	������J�M�V}>��2@$����p;���(ާ�}dｓ�S��+M��k|���&ӂK�;G�����7��{���i[���r\
�DfU�\x�D@�l��MZ���&b�e=��ث�ٱؒ���?4ź��+�b��g��fleX9�����+ؾ��S����ϸ�" "H�1�@�@��+n?W�i���d놦�3�)G*鈐xW����T�?�6�!��:�F#6����q�bd̀*i�T2W�iKPR9Ѳ���X��t��^��p�M�~o��-�H�/�����<<6�=L��������?�pN �]E��XҦkI��,��#�iFڛ[3i�hR}^��D���/�}��J�hw��̲��fI%��f���x]��K{=��K���{�	�S�Sh&b�)GU)˷������}�<���F��tI��?����p�����7R��X9I��Lk;y�ܐa�4"զ�Y�q����da���@�3հ�1���/� Wq[k�.�E>��	�I������*�h�#�mr��ŐtF�����Q���rÏ,to!�#Ƈ�S=�[h������!�:=�o��w,e�5q����rb�E�_"75Ȝ=��w'FBm�O��C=y맫;)پ�CR����Z8��B�&�g�3�Z>�h��Cog��:>d/��H��3�	J�>�ɸ���t�SK�[�g|z<����K�Y�tA�j��FJq&����uPV�Fڅ�D�N�v^�@t��f	.jnL	rf�+�'TxD���g�%�C�S�o���F��6Ѝ�q[3牝 ��6in�d>�0�A`����] �9_�A��[��K��T6u}��{�l�XUT���Zu)-$w��O(�׈�=�'��x��	���};3D�'/}�N3E� ^Oj�LN���#�p��7�$A�j�Y���P��-��_rc�D��i����W����;U/=�y�Vj& ��b�[�7)�p�A��jL.3���c�����/���\`IMv��h_����J���k+��E��ϲ��O.����W4,¢��k��y20�BI�(7�LhLt*��$�~�6�엟����ܸ/Mp���:����w���㼸��%�Gq��;�b�)����M��f�1���ɼX5�Ib�����.�$�s�f�nkL����䭃).��d��/��7���z�Cg��s�"�e���Ĩ�e=�D�/�j���x���R��F)��Cg�*I�ԉ$k� Q;�w[[�ɯy�01�T�#���d��m ���v��0��ym1�(g,˥��t�_��s"��*��q?Y D�����Y�5����'�,i`���۰�j�����Y���9�e9hWFb�aUp w���hF�����j�%@)��"%�&�����E��G0���a>au�Q�dģ���]��\�>��B��`��A�D����_P[�=�ڐ&Z�_J�B��5J�\S(D�U��+����/�&1����3������[vP�D~M����OL/0���0j��?���gÑ�N��MU��4/��8Q=��'U�َ�x?�C�ҁ��Ջ��> +�#�7Z������V�D�_J��7,�3C-pvq��E䵡v��J��DeX���>恼s�w���O �K�����;|X%7_
������;_�)�Lf�!����a=�oR�M�z��ɜ*�Y��n-�����4(/u�(w�l�k��]�n�yjG2I����\�՜l���e�0�{���@$�r��R�$}��J'd�i3�M�,�3����J�Q{�b�U�zYb���<'�ʇ�!Z�AD������[>�9����T���$} i���6"���޳���^�K�^t@԰���]�;ƚqJXvO��_	W3 xQ�
�{U�8f��%TUU$ApgR|�߻2�وm���%�k�H��"Er��u0��bέ*��3]��*Z��z}pS�6?�}p�����l�5>����x�D���^� )�,�{x�uw����i:��Qwt��e�\�K�$�A��pzk�p��y�'����7V:�N����$��,4h�A�o�\ى���gZ7k]�$1��Ӟ�Za�,���s����[{܁�m\�{�%GB#H���g�D	�ƹl��T~���U,;r���S��ԛrE/%&��Ƥ� w��ҏ�Q_�\74���$�� �{Ic�̱�d`�"L?l[�_6���-����mv�����X�V��̈́<�?�ʛ���_��%����t�����-�O�O2���G6�l��bA�ZW5�hM��Q��Z�`h�#�!�k`��kgz�פ�
B=��C@��v�v�y%֐B�%�<��1k���9�!v3� -�P�?iH�����ғ�xa
��`�вȳ�U q�'��:S���V��6�7.��z�+����gL���HZ鞯j�)¦b���ļ�q�Ujԫg��0B����ﮜ]����ixHF޸�+�9�������ħ���?v�b���+�^s���>�4Y5�."��X��B���9f�GL֩���#�˔�ıU�~�ڢϛ�V`�����B��Ӽ�/LO�qI��������=H�G�̏���i�EB!�6�cX���_�%r��Ӯ��V��� �/��C�ܛ���&gf�ʲ�S�C<�Z=:���L� �����h�N��ѠT�H%�N����$ݳ~��>?�k�0�U��PEɾh0�1iP�`b����z)%�Ŝe9��fDV��*<Xc��q�ZG�Z��֤�v̿���M�
5�oh�š������,�>�qɱ�ۚ'������q$��x�+��a���]W躔��f�����o͗� OsS��U�eBW�)i+��K%�׆~��۔�T	ݙ�p�M��#d)�Z�7��$�ѫOm!�{}��:����������h����0��ѽ,������7�H�:�%��O!���)h��(�5����Om\�Q$ЊS�F ��h��a�w�+lۛ�!t+�r
�;ۖ���J��^P�ݵ��Nn�r�*��%Eʗ�԰����M�M��؇:u�o�x�k��-�=W6u��w��r�$�,.�z����-�u9�</HjP��߷��� �+�N��ѵ��X����t��@�O`	|7��"C� �Sbb.n]8E
7���0���=\Y����	i������F�#���(��U#�Kˀ�9��u
A+�N�J����ʯR�fo�a� \P6ݖ���i�����8��^��)��O|���T�wݙ�Jv�ܘT�J�y�'ּ����\1�Ä��b i2��pʚ����9���"}!����2Jz�-w �Sz����,���Y8�y�,�ϳ�y^�
u
�~�
-C*c4��k{G���ɴ���z�c7����<�q��[)l>G#���s�LgF��ZUi�Yķ�	T��~�R���#����ԭ�,�t����Hc`�Uf�e�W���K���l�D�؄�`��R|����>��z�w�}�'��8���kR.�j��6�f�YQ9!��h����l;'"��<�&����S��Hl�CX����J�XK�K�R\�i�H(F�����G�u ~�m��neM�4	%���L���ekPŬg,��b*�֕z����'ݭ�{p���}��	utlY�x:�t!���mI�E6�C66E�W�Έ��"KU��X�>��H�Y��x8��b���
v#�{[��$�>=Q�*����|��i˯��:�o��z�ߓ[��0�~��oޢ���������Ա$2b�p����wI�D�N$B�Ӆ}fln�5�I� O��;�N�jZ~$T�[�Ӕ���N(fOh�{�w��Uo`d�YM�L���P���<qI��s�:�A�������A���4��^�1L��<������b��:����[Ӽ���qj��I������C�s�RW�׵aaJ�k	��gӶ���� .i�O.�rsy�{8�}�{x�t�ԥ���t}T�/P;ǣqP�A����.�R���&�W:[��.!�+!pF�g��K�(�0{)���������c�xUܧp1;isHwc?X�7&�� L_�Ɓ5�鍘��#�u�Ny�l{RޑT�����c,.B�Kd\aXhb8̓*/�ǎg�xQ�X��iq�G�/;����p�ɝ>�8�ca�}<�S]�p:w��A���S�r�� �@�%���z����;��/8�A���%����[Nm]������ ��.y���:,h������Ր����/g�Q��kz��Ug��5ۋQc�'e�� l���/�#��lB��6��MV���yr�a��mX�h�3��G@4�%M@�U����A������|��zzJ_J�~f���$�Q�̡V�髴(�(}��C�׈�d&r~>��ϝQ����|Ӫ�mHFo*~[_` H�r����<��H���5�̭���i=��OG��=~a4ËŔ���UY￧�%v�.3��V+W��}y ��t���ҟ6��Y�2��\�]�dE�ָ��L��"��Mp3��_��Z<hſ��Že��`�vmך�'g�
�������YL�l:�G��t�q�����D{?��~7�Z84��I�yKj�Qi�� ���3Z1y4s�(B��XQj^�oc{9���i�����>p�����p��������J���C��z
 S���h���֬j����B�;R�(Y�h�z��u;}��-\���X	g�t}nMy�#�Kۚ዗���-Ǉ�hTt?�F�K˃NL&3灅M
f��#�);��^tpd�8�!�!�������<���a�����po6�B~�9*�:��ZL;�V�"pm)M�3��8���s�$�ܚ��.���Ut�p���)��UԂ��z�P��.u�N'�~���w�)}�<ҷ�dn�j��W�d|��=������ŭ�M�WFN7)�?9h���3�v���'���^�t9R���Q*L��F����=����U�E+�����_��Od�?F�z�,���]�b��]�&�Xg$���l�Iurߢ�%En4��ѠA�B�����(��+�wIc���x��]��]C2��.�74	�yȕ�mO1e�٣U$���3�l��K͙CO�w(�I'���P��C([��.`���_���l.����!Z4��9�7F�����ʡp�QB&D���'C���(�/h�a8���.d�_�����[�.`��2��ز0�.�=Z]xN��}W�2��s0��u�����<�+/�c�@�r��5��k�����������G�����]y:��x�(��!��c8��n�\;��S����A	�߫��jٜd�h�� �F����0^ݴ�꓋^���i.VYf�5�~��~'�<�mơ��*���6Z����&�z6��zmfJ��[�/�5$�j-�s)<���ҖCQW���Q`:p����)Am�KI�\�R}�BO��RZ�3oκ1e�{��n���	w�uyڛF|PB�Lj�����L�f���Zs�^b*�N��$�tP�w�'��Ԙ0�_KM_���Q�9����~��P�+��h�8��~F7���"�0bY0����ex�
�.��&�蒽dN���^B9��F:Q�����+�Q���1��i�(R*�{!'��L_�ĭ���kQ�Z��B�$�Z$/f�����u/��y�I�u4V
}��\��h��g��}.+��tf(`g���N�|9�t��� d�� �W�-����u��+YW,y��B�z�
��H���#���ϋb+�S]u(�'Ū�0���i�}v_��Ҥ��@�kO�z�|�0`�9�6M�����.hkQ������i���m�#��ͷ+�IF��V�^�C$n�d��Ε����d��BLd�$͊��M
���M�9�I��A���&�J%��81�ElM�	�J��A�cE�4h��Q/�A�W xݶ�9cfL^�y��~���PE߭�A�#�����Ӊ'�q�\A���n�A6��׃��M���/7�zgK��[5����
\H-��G���eD���'.�|=�˙�'�,����6�?@��5$�=`4^Q���8{���c��9rX���óh�G"Ft��H��Y�R�^!Gti;]z�N��͐�+���,�FqUT7�c�1ye�� vy�4h%#y>>ƩZ���~>��#�<'�m����R%�!c!<��d��P�b�qt�3��s���:OB!�j�N���¦R��銪��1�byB��b��2n��A���9b>����ќj�� O_�3��x��0�0D[q�,qNňd��g�u��mP��5�{�H2y��np��!���M�j�o��+L�����VtA;e���Nq4C1�Ŗ�����֎�.�}�J����U7ӽ��F׶�U�a3殟 �C��]<�m�B�@b���+�w��֩�Icب�5D�������Ъ?�Z�H�K3�����8�;�o����@�ì���Z��Z�"�S;Ai���褐rk���Z���+T6�+�B��Q�ne������ꛖ,=�!��q�@g�(ҕ{�%|<�4���Ky��nQg�ME%{7���F`{��F}g��؆Qe�����`��r1�Ѿ^.1(��!pk�0��ʙt>�ߏBo0v���ߣ�/�#��H�eα��P���<9yk,��S`�R��'�E��Ɏ��[嫎!WLӐ��������2�v�8B%� �F�������.f��	���-Jr�_V+w��3�z�>I��R���0�h�@�U��'��|`.��殺�7d��K ��d���-��,�n�3ΐ����s�G�R�ҡ�i`A��X���9����w{�W?|�cǂ`[s�)�6�EeEEq�Q����mb�������׮����U����"O��X-ݘ8 �]��ړ�X��v���ak?����ܳؕM��,Ō`�OB�Q;!F:�$���2
� �g��?::����p���Q{7Ar����� �{9x�\��!��@����$�