-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Kwzxwzs2aV3sqyvnwjPS0MsIdq4b2iWJC9mixr7eql7u9wjMRVkiHlY3aGXdVQEQ059w8afv/8MN
2l0WazNs6D7l9ty5AVxLga3CohqHUIu9qve/RkNi56xLJLsHRO7BxGyUSQvDIG5T6Wej2dwfV0um
oQMKidhTpI9luLcE/xgM0w6CJ4DZM1/kEa/0XGglhxlJpIuEfjdOaB4KcyEmgesfRmVpnjN7hxc4
WUDDocxYQ7TnQrBVyaDiCNVvtY6nI3Euoyo9Hn44UDOlyBaWWo4xdmMXlsdIwA64B07NXVDK+rmD
HBz+TAN50Y8KILzymzZjiJ4L6AoaYo4dmdduAw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12384)
`protect data_block
bLp4/V8i25S9YXRlPe5KmfnYoxU4DHm1u4PQICHIGU+InCF+fVQBIENiR1LYNrnwRhuf9tR9cCG4
e7AE7K9hinZSvp7xFTfNkO2/qksGU36Ej4mb/gvqwYWehrY/XGl/+KOvt30mJ2wi70CSLSJqo8R2
rNdyGdeOwWFbgzlNgFTtccqOx1YuxNA3VnihrpC1k36PM11gSHVGR7SrHGMeLEH5dKOQJaj270J5
Z/m8wpSaf9SS81HXEuOxpKe5nBP4jSbTwPYZyRe5319djkG6sNZsv76GNLDQTWfYekCvNgQZ7v3n
u2xcG8uHJOuyUQtGMmk7/BxIHiyhthfavolzSapXidEi52Sb6LrahGK2zGrgvS/X3/uo00Cm6Azp
v3JlQQH12U4N6SMX2ZE1zq3cwcD49jcPrcup468kGgVZzzNPdUnJ1d70JBTrNnN487g3FlM0iOr9
T5Szy4wpH7I3kshTQSYmM/d1dMfKk/B6L/gm1A9DSQW0TvPP0Ys3jB46A/jpOJvTPU8VgKDliGVG
jYWbpu1KuwX5PL5W7DKTZf9j2z8TFOtmOfzC436IL5ShQDYUDNvJKA28HOugPaXmcju5ndivAk67
uf5pS7OPlBK7dKaHeI0wLm3fGKvPfPh6mus5/4nmjfTfwnJkRvaTkKI6AFmqnHpGF5NNCwL6/G0J
mEXC+rcsRN0yjRGAAIKwWO8pU63wWJ7lyxs94qKYbFO5za0Zay6jfs76CYFmpSD1ucFIrZkSihpC
bdfzoTDCYFqdpPBlHkPexp7pyQJWnzELYaoB4GVtFNkuoocbfJcmrY2qwtjwU7uTyyVln6VIVuGz
UAihKsW2OkRes7IYclB6F8Zwvbq7undcUAK6dZrhF256RPp0CDEGjB79chBHxbRBwhSrLFumk7jN
d0fpRU0oOK3eXc67pc5bWP8j8a/lyBzUA5gwPJNFleb+6fu1fbpVKhWjGNXQX6vbY8sxh3WyoQIY
I9n7OcPlq4ZFPrY/nVq2/63HS0Ow5y7eMaT/Q5BSzkjZB5Rj9p6F3Yc2pkwNtMXwAC7WnF9X3kBb
SHLkhhfSSbgg+3+lWVFsKf01WHc95wK30d/T0YbcZeH3+vx7BB3oMIYtXpHMhSnQfHl07PROWKm8
Q/qetokbZxmMkVNClY9T6TBC17DkJmCVX3jmIzwMioq9pYzHXOYdFmMl5bnrrqdc+54PraAcJY4O
GgRyVuvzojQTAw1efPW4l0nagHeeSrB4AX73CyApeEZAEzqH76BNwZlqCMeXUC4dOZEgPUIE1n64
as4219l+q0uuoequruNIBeJuTjm8uGz5dtSK/PnzV0cANd/u1INcScVb257WNBftZl+QVLM/4JGf
vnk3jQDzq0cyMMue2mQ1hnqrV0ycyCWnEFswPZKRim8Dv8AAMl3b53tQzj9en1SQVDcneQAjlYO9
27Qlp26WIEtwoG1IU1StLy6Gs9BKSxFhVgfpdZmtce/4NV/3YzPkOcZqW5yj3ZNrrG3ey19UBY80
Vz9BapJh4CQI2zWXt9/iQytRjXXrlpFufG/DDAG8TBr9Uz7/QskczR4yTQ0PZrCuBu1XzVbtGAqg
xcn+IV5UzOREltY9Bjhz4lqfOPuWhDykLh3ISextaxQN8fJeBgrTjmEyxB43XAAFxWU0CrWxKirT
VX62rIWyJHUsCYG7LW4VG90lrfv5rDZvEMI6XDkc6LOYD7XrxoIU+/ceY0+5rrvVJoSv4GAV0wRf
IFIsQef7Bxd8BVZb3ihnNj3etRbvGweYZ0yHer3V9wo/Vw58mSBIleTywTlt0A0oBld4+0YnBphQ
BGUexCdm79BR6GZlSJ/Wn7wpvgYMpLwM7GOqO+Z3g2nfEnM2I1KRPxSVWjhqX7c4tK9v0MfEwUCp
GQkLKTC6BGJIUtF4PC3kbtWy40qtW0VAhmLuKALke+LWm8aLgkKL8A52Yl3NLAtx2e63xcl2tNq1
i0aT3MD9D3LnT8UfYodOFyn3GFwPuJZ3G9Uxo9KTR0eNhiXd844J6YFrPaI0kJRpeQ97qkDTF5Bg
ModLHfOoOhEPiGFSPmiBz1RN+SXqL3LlQZNH9SDAnMp7U/zoUSLxDH43jT+WPdPYJygFo+XaDKhJ
AhNLMniJJbzveY7xeQHTmO+wNysapfRDyT/FZpSV7OSZnb183BKRXjxdOKehyWAlFRAr0yk2Drjd
UQoX5s5d1+qbctMhDd9njSuvdOWpLOOkMdfMxFW+xzBMK0SHqbhgY6zaeMmpfVKUP5/qp8iBQAUp
JvSTzfsdO628hcbDezxDTO47L/C0QbX1UEqE+yGx+Jvpxp+SBwukoXAG9icVaK/4BvkRLjDgnAcc
2wHNq9MBjJg9H+sDqXrdxPbi+NdKiwRDwoaqiZ2+ZN69XuHzaM7cE0fG8Wj4fJGUOXRO3++uzwBr
OVR5l80qmlgwhC+Xv9K+ePNEed18kcmEqKE+Hfi8wQW5YFFu7g49HJscgq1VivhdkgmuwjxW8eUk
lD/rFz0Xft6VHE43GxwgVLC3UQE71tICSeCF8JvCaHrmR/r2xisQFNcKimGWd0gS5UCiZOxQsggg
BBeFXYkKxbb0Z/k/QmeupwrrNG0LSu81E3+M70yu2q/lbRHUF50FrgeN9GyNnlxuVnsLy2dSOY7S
Vm8JqQX/Yj3cxLMS9UlakVQ4tpqRwfEuDCJyBl8v3p8YTZMzTiICmGe+YECdi5nSx3g+JdqENd+b
L7XMEFDQLY4bgCLy1jULKTAZzqrc5LEGu0WCkKbVK9TvjMeolFvZSWgQtU4SBFDd/NYnBkrrEbUY
fVbUcc3T88WLfytHjbUFks3WzJHjvP4Xq549yHBhvoQB3k1JIbD4PqDBPeNNsN2hKePNgpNaJhhg
TzQ0rrv+Eld/K0Z/AAq1nc/yPJx3U2h/3hwy8HYTqSavlzTu8/WGR9mROei1B50cVQKEzQNab1Yk
o6rLsOp4T/evwG4j7di8ADItPfNIjwMf9efEOYyc9hDml4Waf4OJCO2dQXV1Fp9sXy5rwaW1lGoZ
eyWPZRfmpEzCMCJlR3Ovsu6Xd0bHG24PCNsgt8OfFEjdWSfEarIyvtcMA0615JRinr5Bn1c6xRbe
LAk8VP9uxniOXM090Kjf+/O/aNfBz4PpplHjAmRic+yyIp3tXtvm3Se44kbBoth+LZhNNXin+t76
OBGQbbinYjf9EnwVcREstl7Tl3+P6YABLVJGYRLqGPAvd7dEQo8gtdXmdYCFVn7XxEpw+TxNkOb3
UetmwvVpDouQaQlVch72Peca6vnSqgqi+Xjxm0oxJbKaXx9ms5CyNfn3Fz2PUhLVy/hPQ83D3UbX
4frTEQkH2YcU2LBy3gazKDO5pL8iitsgkRJl1V0l4ectPheq+2wwGZHYERscy/AZMHBbt8IJgeIh
CxVC+nJV7jsHcilFqcY3zcMrp2oSMIkAhtl7jpGl8TiTxouulfWG/HSybx9WZtYf5hsbWlvyvRZQ
R7RJ7xzZzxsqn8csY6zW+gkZn92/3CL9aLdgfJEIUSJ47+4A2F4ao5/gH8YatfYl6dk6kFUv1uxw
eOpYdsyqofjXH3AODJ3mgJ8VoRL+z0PPizGMnQ32AmlPp4IKHQA8d9xpk6swlZ/T4Q6z9BrMlO3Q
BAUJ8o+EOcyunZNQCv2boV4O9L1lG49yrtuNzWPjE1B0lNIKCEMSJFSadY0WJvyswCSC4ULPDh3I
nNnuY6adFaRmu4W7EBEx7LgGDwExYA+n9CRqA9sII9k04Un3u22zWvAF6fElJOC3lapu1dAODZ9f
RRwSOWAaNA22A2Ksdec1jlAkkp7cOqburk3xiWoRyGzOOcwdyuAUgtTuToQaaYD6Iar1B7UwkJFc
PfykQcO/RRuK2a1+onTMCv+X6FNfV7PVt530S5otDD12mN0t/qbihd7HM9HUAEiXVXX/emJa1fE3
QGSIczWymXzJbdSPm+oMCtYlBOrLqD4WvSnXp7umqKJpwo73iaLyiF6FD3YoNZUXVXo0dE7omU31
PIcmRZgQQs3a/xdTgb2zdHb8azHhNICd0Xe15MlFPi2WUbLkxIA+j2YP7R1Gfa6LznvdLqQ+GxDp
i+ZN4S1k+WD2HjwDfBn4ubAT5pPVE3CoM+5hn+hY7hsviK1gb2ETIAwM43tyBG4csBxT3ODgF8FN
KEmjxrGQnKV9Try3ySo0jLfE0pT84VocWyDnEP/PvytgvervHBI2grXAkWLamfvjZetNmp7AVXWb
2qH1uoQatw4zmjc6VDZYtZt+pH5vi/1g0Ra8Dpw1s/LFn0x94FxhUdnDuKl1SG2kuHuJ0HfZuFdj
2fwGtOvECmcsDSFCl6Er/gUK8Ac+qHFYuw3K662GYe2rIfJOhuMEIrJZuaIIVPHly4B3sA3qpAbE
aLM36d+Tb+L6Hv9YEUSOWZhgCK7CSGfvNTxpQw593imrdBmqIVF3ETMcz09SVYP3Yn0FZLO1Si0n
vYBstBuqdwSoWGnDEqsuTEGifQy7KnKBJojyvgEMJG3mcWfwhgWLtVhzVhaYAi632Np+1jJn0x6H
TTtODRwuuMBu6a99d0ykzlqPyQYrlKp2cOq0aElq62kpPrY1pP+dwG242ZFLd//wVq4wP70pga83
88xD4yyu0GTS86/jeixpaJiGySlF028qJ1Nu2UfYVJ91QX78FnY2ZZiTHhRWMiv9fdKHB1xqO/3w
pCGf0pGuCmLA8Zv2EQd99m5+Tl8ksKbWw26Xlfo+beaLf3X8KZsfGI0Yvzt8TdjcPa0IevaHjACO
zCaQB9hGzpS7MoxQoi/n3E8hxKtZ83t4weUUwJeEqex3mVbsa88Pd5nj1r7ANwWbWUSV81BksjBL
sUeAv2M9g/E6EsqZQrHDFrHDM2UEujwCEXK922r+x/Yn3+xVi6BOJfV1DxIMxyRVnBjKW7BTnbaq
fR6t4nkEWIzJjO/WI/YtA1LvoBH1G3Knf5L5aB2KaI7ucGeM1UAbTTbeSwkfTrqtHarh2V5dBoxq
fr0JlGSg3P+0XWEPq8+Ev8YukQ0JLEXDTglf6wA4rchKiS21i1dXy3n3fTt0RXbQkqR28xG9KjE2
Q/0wcCtIm7gZByPMtfPjqfA72SFYv0S6Dn89ROBlvSeICsRzv51+SwoRh17SG1P7YIpZ+5kxslVb
EUv6Ib5J98fSLTXXHygev4XE/DbTKK6P9DJiyqYwrM9sxPR1syzWCpV6EvQendF2ypt651fN4DCP
CRcvAlw7QxAueNoqkeCiNkgpHzolwDvqsjh9n9jXceon3v3gv+c4cFXar729DQSX15SoywHV4spN
FWVqI63Y+t68jNBRvFpjrnFqIOaUvthLtc65gNWykB0qPYw3Xog2rktLEz89AU1nENhRMYsaC1B3
V5+jf56NdeDfInF1yDCLBq6d43iC2A1rY8tULJR1JkxLG7PSJbpZnEHcZA6P0andeXEUzczOcPgI
NN1O4rVNpvcRZUDi8RPbCdSsWyncLtGE+wJbm2tcWpEBQ+9yQxYJJRFCiAgaOXYHXpiJ/rD/AITO
Sxa/fJDLvgzkwApCwrxr7KW45Vweh7HgnSGnt4iqbia7hGZbABKrCYqiE4HCv1q6dAXHEkCjJ/uW
4JiK4WEbdzkkXXpocxHeGLasgsYvCmMg1KeOI/JxW4+5hSGbV8zOjzKBiIbyrpHjSdfrZxKmFKrV
Yi5xVvwCSpsWr1FwTbeNM5KtZmtBCwTjHqejgSyLP4kRgxQ9ONuwzwpuLiBB9AJLdhfSy7aMtaOL
JBeJk7gMZ+REmpkNXMPjJxuvTVRxMjG8hJQszeVz7SuVsS7j9Q0Ha7t/MFn9ycWBTQIHvwHj5z5I
ROwKHlLRI+aalxkMTakCRUD9r4Nt3S0jOY9wOXLavmzq9WxX+1QzlprEtEXgAykjjEdXH1afhqGa
k20T729/+QS1whaGxGF3Jf4MtoMNERheoKeyQIZW3PDunr+5fj6Ux9Qgf4/ni0cNbKYIqxo18b2k
0JKF680QNLdGcHBLLeShPYOcQfyWNrAqtK2LLE114x/Rt95LzG0dpVCTLvkdrvOtl118Eaw2aFEs
SItMgHSE36ETP96SKFJfo2WYi3l52IWSz3h3Fcxikae3l8+xXv4iD3hMuiY+ZxJsZN8c3xReV1tv
r6vv3CIrXAzWXLLCaeGBS+7HT6Hsp5QVfROjKRcR6HaMRuTI6LmmeogYw+VAHVxg4YzwcxMnY2n3
d2ft4WxpN+QxOepRnU8BTHPbfSIYxHk7EB5lRuBOkkFy6zYB/iQtoFSAkg2VaG9ZgMEPdnXJIp/m
3UTIw8oj1KjC8fwIqsDBIa+VJRLUyrbfwhixz6pZyP4SNoO4yjtGss3NPQghMWa2TqZFcejJZxS9
R9V8wtOquKcPKrmXOdqdq6xlXyYeOd4SjOLHtK2qTtrHT1HVmVL0rBA8ZYyjmeToMJ2jWaaAeBcV
BHmfklR1IAjOA2nyGyoWpjEH8YGbWZ6dBpOMDOX2yIdFuIBWOEnaMMlZwu0X+R1XdEO9CIxKRYa+
jnGdGo9hj6l/KAtqE5XZ2WKukAHoPrsEXI45EBP2Zm1A9a4oy+1s+wIVwVt8LcXGyUZtCZcKtEN9
KKVkzQECDhg8Ecp2Ay0+YfM5lvA/UfCIzfsfqMZjQ+QTAvnoiHQjG++WRW8rt1uA+H4KKH2r5LOe
dEaimt3CbnydXv7O3szNkNYE1LKyq3Gv+wmBGfW8C/+hUgt+LpeWSOBmzukLTDXc91EGeNOwgFVZ
FbddRTISHtS2/KRvKnaCGrAy0uGa4HIvM1eDx42uitszLh8WFWvI4RJ/w++jsg4rrr+3+8hW+1fy
xFdIwkliGkrjpaBZRdEZPnCKS0Kx6ZkYsTN8y+uL30cNvjb13fVPgS7MYA6VLlIM+cnlWi7ap2tX
bMN9TA76IRjqHOe9g64JBmk5w62C5hNU80QZacIZJNQL0q7I7nlk+BMzVTAo3wEtfCMSoShClvNM
9cwu5lhu/CPM88MEB89PSU0EowWVgAq97Apf+nEAvE5f73Zphb7dPW2Q3uLXYG5+XP0PffuB726Z
eMnnlMNga2/QbHBOvHT6GdwmuxPStGjTQXQ6twK1XP9aXksjAS9GOoVb/hGQGE6BfbFfrfCiz34E
mb4XIkLtSX5Olf5lPkD05dA/Hv2ev/Oydo3/Ehai6dxNWv+z7Bwodh+tLZH/Li6jbvBdEJQ/1Ff2
TQkG+u2SN6rOql+wMldzLQQ0Ea0vrSNVQf7Q1dBgrcggbNaeVjQIsbMgQd3QKABXMrE0GB/MSoJu
ncX68UI43vmYML2N5sIB7Fbt+2dAhkSlTkIL4iNI/uOk95WpRXyYAANMN4pbteEPwvcDXYayS9+q
tbY9uib5267FRhMSORgXm+RiDP0zDXFBMVXGqd8ur1sq7rglfbJqMalLml00KvRyhbp3INJGrqJY
6x+jhqFclebwXoI6ogZ6KfXWFijYFvQehedCW+E/iHQSIZD6h6DN0ODxr1MGflC8XX0CGPDk846i
0lIcTNxtoc/mc7xf5J+tN62nA5gELQS1EkMSnpa6x8hM9Dh8wUcJVtBs5Z6mtnf5yy0pmC3rSGXz
W3dCMUZESujjMu/ZkzFGVOw1nnzDxnPzqogdV9+kSb9iGKcxIeWPxOqN2PIgz0VhP90eUVTzcCq4
uVms5q/iucfWfKmHkzbDt1ct+Zuyn+HrcfP92MQhpxPeoixmBx/frLnNfyO5XI4tEZkil2W9f0Zc
ZRZapjhpg6OLh9WtYQsT438/k6aoaP2BLHrvZJhOZ1SplLgCM2Qr4shu5xHDqHFLz8/Yum43wSBN
aGtFp5F5sY8IY6RuANnNXDa2NpCvT44artc00xukuOcuuCqcXhNhcRvfwzRrvOY4DXv1GSB7mWHz
WtvzMe4ZeuLLxL6j1mLeBU3BGRNWstiSC12yOjtDn26V8uBgkGeYPMx270BF4es+BIjYIYalmzGR
8q84bB+k9ENI/29/fxXJ/ATLc9yT4KA/KmMwefzWD16sRvPNmH/aKtucic+k5UaXqOwKZEjvkuwQ
Y25FJmrLZRrGe3on9Se558VD3EUsTbPGsCK0Ivo+qmAUZyV5U4NzCuUpJh7bmpHO7fAhyoyt4SeO
3ih59LcS6JtuPitHHs38XtTrh5FU0q/p3Tc1TvSVuGeeuS+uI/zMYkDl7PzmwSTweU9tuFnkIu59
PHFWyKZzO07+SB+rQ58AauNPXV08JQM6CP/oauroVOIvPgUwipKHPGh6bmT2ygEmqYO62jU1ENU6
x92IiMWlyG1dHjih7pRsNbz1tqnN550Q85Lb5dHsLG/G1YVLmWR7l9RVENEiR10yAdIK064itN/N
U56eie6y9FNJKP0jS9aqpPQhFimOl9Iw1iSXZvO3ODGS70BfznjXkKErglKQ6C5UKWmmfxj8ygVd
ZpdyEmp/Dep5yFxv1rni+8ns5vCpd0bcUnPff1B9nVTQr+xYBUHOPnlFpMdasHyUG3gL31YEY2Q9
PaSKxVH1gcRjVR2xKBAv1RVI2lH7Lz1LJTKC/vo5guLQBR6V5DIPqGFsO2k3ssBXgXTNAo3L77Cz
PcsijIcG+YiKJQTZ8+NJpq9nJ6UP4ibAzLGx4Hx6Vx/TorUMscGF0FozwCf82xDOAKX+TORd93EO
Yr10PsXv/14PSv3HRslLFVl8LEDdz74RDnIUTsb6tOcMVKNz9nirAD7VUWj3CotTMYYk0IcTly1u
GYidYRRTMH4JImSE0Fa2JcZLfoJ03J+BLx57jJBBjF4o67cLCMuK+WNAkgrrKSlA3/pvtx1Ybgem
dM7W+/sJQ5WOH+RwbATQP48TabeXBGrOCyCrjBAZKs7Atn/jnA8cT2WSzfWoLh+IPWsXeoqoowrm
hs3lr2do4QYdMn5OD8CFnRnGcF6lGNTj2WCVkV2e8hXNCZ6cGLa3ZVLokMJyFp/8gz9impt+Rcj2
p1sFpynqPE3uj/POUd55b9oi8naQ0UYqtj5QOr2589fR+Dcdpudhn/ECmlEnPvgLoH+VbbrdSk7r
oBECBbALs533QzuzaJvy6VmLLc1jtmYnXz5W/BARUBL+Wkjj9lbBEoObYvKYcE+CkoF5YMfLlYRm
puH1XQRhJm5VkV+YCSPNCMrW4mn2uJRRmdleL3lho3qsr3Kuevbjud457XSTdoe2MlVg07lV0gDa
9J9b4mu0Wek+7fWB3XvN4DShn8C5RGRJSaN7rfvIrLSyS7XZa5YPLWXgfexdX7hQ9zYVwSZ36Dlx
owMj9EiDlgiWbl2a0Tdi3pW8j65c/pOIhNPerOoq1GTZ1QJcYeA3LO5obSGB40jzr2i2fv24s2gl
edHLKqraVGh7Mn7IZ85py1IZyUNb8IvSZBHziAvej9RplelDiggFYpPnau0eSl9aWxO4/zWypGG3
UvxOUZCTMVwun/0t9hC4Ofj8IkPpdfM7QGDI9KMXhBzS8s8EwwbO/faAtu7a5Zk/Z6JScHRQtFI4
aEDXD7Ip9b7+gVKGwa3/QiN71wegUeSXyxLI17QDLe0yvQL/X3wwOBWNKvkSnGKIMzdPFQlp57If
2hgqUCNViig69AnjXdWvd1v1SXDWsmUSUk7B3W9Qifd22oatUjWwRjld4bqKVKwgm4wTD5wAOVXd
+EnsIIXsDCgYgHo5rSHziSwWtnnC0sddlOEwuuAr5cC+cFkQVrqqgQBp3Ege5rqK3P5+00IRt987
3+/JLd2qgPYpZL1br72oZl4wjY7kQti9PyY+Nk+lzLNlXXW5O1CB08dGeDI366bCDI8ZeJ1Hsyi5
326PDcpOm23uSzrklmj6roQULbypP+Q3vCSPXVxQ1HPvkjKUOrL3AKQJQqTV6d76VDlWeP28Dcws
/kXxgYcl+3Wj41yyPMaxZ0pJUxG5A69t1/Oi82ci1W7ej+zt1OWl3IdqA/3K7BVs/qIRK8lyAZUh
45jtviJ2RWqCytep1dApPHWQ+Anzx8USdnjtCp+60V5/rA5XNe+UJ+hlxw+zSm8GHPvo2GO1AsXu
RYnZOS0skk9jdBrWX63SQRhSaw2AD+q+fNVJz2nF9XtQJ/AilVC5KA0nc+15fa3zujRXm6wX4I6a
RZ7jaFO43q7qVJUyIz7LQl5LgZgXxamOUAXydMIf+N0PCSIOU2ACB9tcNqbOfWxZDDvGv6fQIZgH
RyUtDBSkrC1wbzOZUwxfTOUBRzrXMxOd2YgVt50hZU13mQD/Q/YXqM2nzdoVMRVQeqQ5mghRxxXZ
CI1zWLeW5ZhvppPxElxdY9TaI/VpXgBfmP93YUFh7h14VzkkEXJca4E63ML2cXS7/zm/gZ499HFh
uaKt3uN5fg2UpfM5prd7oPZpgAD/9wDZdz8GLXjr2VTmDoHMZljoSq7KjwoCQwEgsWAcgU188IiJ
9ms3Yi/AskY2fPsHy10I6nFWpnjI19aqMQ8XumTXSICUoF2VRwUQ2SizGsnox9mEyMv2dEMY6rXq
CNTspAjoefafYawkm/KFQi8auHEtUIf8RTnyGtL/x/l+CZwGpp2F4mERDg4YtmVFYTIbKqNT+wqh
W2jDPby2cFOCtzfaOvkVT2fbvwBKwZrU3S1UuPYwnm7cBGsujafRe8DkevMulbGAuzbgcDjRwN65
XlxZO5K1QMfK90mzql4hpCZRB1Q8Ai1cshY3DTZjo/s50s4IFer8OXywMjgdzDEn3PC++Ems9i8a
EDhUPxB9SW6rskjVoxk9AZCPmbwuNrrojfn5YBur4seEsOiRCIjQcIwTbCitPrRxqw7teM721XSg
QpS3ItwFHpiQ9JCVPgeWB4uhpQj/8ghy+jfZMZjllmLg933Mw/4bZzPtW2EWQDRnRzGqDS9lvPnt
Ld8pcy3n26M9UGB9dsAIGGqkRiM15L92Uw+jjLFKaJdrrRt1hi+eNdzf8/yvVY+JWOIyooXHOFSs
JCbPDRNxBHfK+p2nD/MKDUsPl9jO1RJXIRev5xM8QH9bGJufreEGAk9oAI4ZPXj1J6WoVnoACpgG
jx2yrEcjAql1Tf2UWtjFkpBxOI/yRnLGEbCVwsHSFPKnVfCvAKVnSus9vuDobc/nuUt9U3nhmAey
8ludpH9UpkVEpRmrHLCscO/1QWWg1kTB7NICX+27+G1c3o9qQTX4XmOzxYBUvTDmfvJQN1wFDHtu
F2R4B3YrLfIhDevg001evBXgyrYjJrzwBlCukbTGxB9uvPvocXtiC5krI8K9ipwBHybtF9tK8fWt
B6Op3A1y01VD9QoyeQQ7QStHCNmW1b1FZBIe775svpWuumd6DdatyMp29zzps25iSTpTfZWEQeIU
1HGm9AbNtyeOCFKg4tJzKy1D+SkYss12vr3n+gXnqU0Nm+KWXg5ms9MI74J0JGr0IathTzCGpYC4
nfWtX1Tmj7dAga+JWAkuDzkRTUUIgFh8B1cZzMS4+fLaZb3vg8BXCm2mC0rpuzKYr7ubJ+41EMeR
fuqxS7GZgYXNKBZy5sSPujFgUX7GU5QKLsHtH/TvAPB/qFR4VTXVt1h/O0xYZYI/4/HrBGfYAy3t
EXvGsWgLj6mUr9PJBUG5Gc0X+QLy731iOBXgw1ipflSDOnXRvGUvB+YhVvlxoomheeQVmq16zDud
mTDM/X8jKNlTCXr4OfnJ7OiFLm0ZXep1SQE4z8LcEDCdvNG/NTcGsZ9SPOjznzMHD8coJP5YFWC0
0LUBvonSwrciUP78EmNEyzBqSFStGRjFeXacXyaGLu5TLX30j7Z2qqx83feSQS/kFaXx81FvDks2
hLC40vDgTVHn3/53G7UZAI9PUHzj+hYK1gtKKkQ+JC3OyXnb3L8a8UCGmtCTSYAqfRpqL7hC3F2L
K/yb1t6fZsuKbCZU2xwBKN8t9jSoM1R3/NOAC9fzZRGoU24HXsq2/oI9XUklbXFTILRjXawqxz6E
f8NzzyBRwXcYxgL3OiykHQGv4MS5XqHHZsK3dj4cf3CyESlSgL0NjNSdlte+hkrgsEtZbSaJqr1Y
7exX2WEe5q02/U25ddY191rtW/pPV8EGgxivWHGQx26P4dgr8ksRuJTvO9RqMaltQG8Y2jdCsewM
Gjwtc+RnBLzy67laUsohz6GEAaQk/5QoWW094AEALOJ0qndtaWPxOCuleyvxSBkMYnbpEEeIg5ny
T6nNt/OHgVnsmqS8RYPgo6XsF/amtZPY2wNtiDamCacdI2eETtluRjRDIKhFgPMtOkHlxUj7IwuG
dxVQqkj0x+IBXXUeTfuswXap0XIYZ6/44/043S+z0WcPgICbvpAo3D2Av9J+bcwBPhz151e5sznK
SQBWWQBj1l6TG+JSyTy1xHal3cIS/f2Uep5/NP+t2UFNKCcad1SJnljujMCjbBTaDvicswzdG+Kc
+i7xp4jbYMnyx0PuHt3A3YAcVI2B9jftlzxpCUT+ir61Xhd2eoBZkeYv64RbakqC4ZwuGn9WeWzD
fnyizRm9iKlAHfFT0KIk846FPi3P3my134OFYrurnwSdQ4Jgycv+WCj45LGjpxAycr1omzmTY0wV
SpypjxpFIsKYnQAKU3s6H990RWxKBOpOz4z8GkEIe3iLzjeuMBPaAd8QVryVVYv+7sBAK229ylNN
H3idPDRfT773PW8kAfk8SGkrqRkneuiDn4R/ZEM9nY1fVad1sFiQR8MSa72GAO0P2t9JJWq7m0sS
QJxOOscl9MaIFsxtHQ15OGB/ZQYxYZtYI+WfIOlYCOFHbAtW48MjQ/urXlDY1pd/uQVh1PCSJQkR
GQJhDvDme4+0XpFTbAvogmOfHSYl13TBMrVyiTxebJsT3oq3cqNYd4BotwBX6EAiNfYEFTiIFsAy
6+h7Z7PiFw7EIvdjz2cBTV7wr0haDUWWZJf5pX0/po8iiCZfqjmwMTxmHT+/Uh6ZvNKeaaV97T6B
W1rJg5N2oKV5/6/LzhMC1oGsimyOEjiOxjDftbk2urqYK4aqaIU2XshKeRzoB9QoIpgAEqIYDlUe
E08Gtd8BO8H2Kq+sF/WAwBnPvK5GVqPaUwJawEF1Bab1rjL9bIEmK2HVkTZdLqp6o9MoM9PH8dK3
BFjXixdR1bQEyAyPCwO7rygX8vTY2gjueIB2i6DJWv9T7YUElGi12RvwzrlhTx6IQd+ug5J5CnBB
lUBw9+kk1RwdPMUIQSJ7FN4+Xwk1v65iTJPhPqHx0k4Nw0cDIBhlhz91mgBxfeFWBbhk4bQraKaS
sZRloOSL8RXHE6yCXej+/xWKN++HPNKY5Z2PFl4gM7ktXt8yrqq0xsfmskNnTObWkgof0bPVGEC7
U/54z6b1pR/LDDSn5XAiRqtBjzY6mk0wMhjGDYY3dkxL0NQT/E57mBsM7dhLEjcKHC2IMK67mHRr
fCvOdbPj9CNH4RPuPRp2QgU1FPSlevvI9cfg36Mz0O0EaAVHrzQjngL4xNjd0xGvx3grAax07Jsk
Yv1vEowUwXkhoOAA2xUg0VFfmA9qn+KFiYjIySmoVNTZh9PLcGehLNESz0mWgu2RnG6kgrWIfXh/
81MtwQQTAG/iCpZ0SG8+UhtDdEwsyBjqL4wPc7KqtVXe34fvh5FuWJPiVK5mrgI5OY4svmePb0JD
hwfIEAl8Mb73qLSRWnJeF7zM8aM16hxnxCuzyUkuZo7h1MgNq4B4kZfuLUErt3Upa2IIutbomBMM
4/1Olzz1iO4Fi9bbekDdJD+HXuDGgaVj4jfztGWtujcDgREaX6LraBbQi2f33gvb6gHTpMRcGEtE
snsCC3cmOqI79/+Vwko7o8eWWjuw8QZfFMt+Dp2xnU06EqxQ2qmiGNTaWCUkpJ091991y2afjJav
uddTkQ1l1yIqr7FcaySSFarRzdfiuTtiF2UOGmNWA2tH2R4MM4GBXY7bCQt3D91lDBHtQEpICWEq
zckmItzo1S8kvfLTNIQia2oeoVkrePajik5MSXdBzL3FWBNtwexAaKrIz6rzJcK5yn2NFeyvvQUv
z7YstU/Ir3OLYczegQa8LhdTcjqoNjH23KmfxOO287+/K1RVyGv2gJs01oL3E/VFHFg/ORYEHkrL
2mt1OV7g8bfeGxFTd456IugtAnVTuSbIjbu8O2IhbH3hG5b3BJ19vgUaRI4uMxZ0XqB/uiVMZfCV
4A2O+RWRXnDbFs3sP2pqKCMwk2IcDU1uuNsjcNDkE/ItIGxcsl0+IBQrxVH/MNOnV+4z0c/pR9Ck
q4hcavUw9SHyYRsZYWEcEQS6w4ymD1VDum0Sftfru8Wg6gJ9uFQXFwLa99xRje/k0GNbjwlNplmn
WUEHyimOofKe3L5B4msSeCXKZsW0R6k3hMvDg4OPiry080fM/pUAS6Q6Ca1iGb0ptnDWtvCh6beM
7bMDq7ZsYm0ilznRW3F1F1BKKtyF68yiusT3e1GHWxztlHhH5j8j4FdpdWn1CHALKCtRXDgTbzoC
r/v31brFSq8o07E2S3yuRLYfUTRPOzljBo0l8JfLJ5mmAIkMARpklPveINJzKCDMWuU4W5RE8Iq+
Hb+msCHwqt69Lf0E+E3fDtE0Asu53ez2z2WQzt3gvoupLd4tNqsuICgGPHj+Sj+ADd1EV19T8L4T
CVccTXgOHTEatK8FkijIOcAkhVMm87eTyIG5mKX2J8Un/14hRE/o4ThIuvgBvOU4GBqv2L3V9jHq
b6chWf3MzR044GnZDwKvVMhzbAxlKk/AlSUggFqPFd7zeTf60f+zg26UMBr5Jj6Xjn/rVvWNQhRN
m5zY+ia1n0rssz0J7NW1OiFIThrlAORyxvRLRhWoFXpl4xxaMl8ExWAdEsYN08MIQcD5ZtWqI43x
ZSYc6FUNUYxG6aygYvcjEJ+2OhDP/6hP37qWzmkLe6oyNOf1YRdzjAI27EE3MDIEj5qrd36+5xXC
gd1bxXFpOZX8j/ykw9zmN5VINuR22pvOsnqId+y6xmMX9ineIq5TdWNlXK0jh5iqRl9tIAZMRfSF
LrwMqI3RTxjT8yK+IAVg8YjQUYe0vx/sMPe2EpHzkLuJvq/HKT6ixRX/rODuYLPdqhTOtWw4ukOL
5AF7c7AK2DEBjPyUTpB9R6ImjD9w9/ijTATFJEFpHzjtCb3RNvHtMT28PloKCLBrembGl0gS7fQw
Qoyi2Ii0zKK+geaxGBZDNMAnLKRodcFzil1bmd/IEf2jzQtwyv6XVF6tSf687/vq3mMZQGaazQ+n
hzAHbr/Tp2GqfNYWDjFbpR/uSCSaQ7llQoyazl0hqR0Xs2IQMIDeWcngvp3W/C+jWKdGyeYEG9y7
UBTGvBUInF21bTY3fUKzrfjfsksY0xPO8DeoUt/S26xlrudla6r1VQc8oFiBzAVd3sch600xXNO6
t18IJBCJSTXE+uWWXvg9RSHzymn9llH5H6Bg1Kby6iC4cxiZztWqBxBZqFvg6J8DciSLql64+F8i
AMO4eDQj/g9iQ1MKpEzkbRgCdAygppgTKJGr3x71TcIwkGoLEI45xfCEBe/pXf+ea5QqbZHobzlM
+mrf6cLGBnCbIa6WmslCpxYNhWYiPikjiu2WqLJteM1/FsbWR6eyW2+ggGumcszvv3j7W316G2IX
dxblmsneRMpleGeE2lgxGgawYJAouLDlkDj9CXTstcjJVVy6Z4hibTXWI9rdi+jvtt3WVgRb1PF1
0QtDUJLodWHtIifVzPG1ydL45MludEoBHUYex6PfS5y03kphlGdC45bmCo6zK0W2BHiTJSqQagDr
7t6T3eHm+le1zjN/3rQsXHbgBEzxtdycoHDzxwdZ14gSp9jOWbHOZIzr3wo7HD09SX1uv4tjLiEs
rNJ6SVgVVSxNezdIVF/2k00KLYGA/ifgdD8Jcfjfz1AEfb8PoZ1xQLKaan1sCCxMYCMAxDFdtk9Q
PHnk/gnBv6TU8CpD+xcZukLoY3RXAvRjvX5C6N/zVr7qB7fWCxuX1/uES4l3IT1Cyi4FHDo06Zj4
YaXKlhGdKBclKMzyXC7X9noWcMrUNLr/2gx/2FqgINVV352VMCnl4DIsv6eOgZB1gTFL3RNnKd6p
QMulLCTfOIJLfSznQGzdgvoHQUdNoqeUsDeJ/6SKL+enkYQrhMnhU7hek2DpydaWA17kZaQLoWLS
qrzdETQwxrOTiT4ip5NhpqkVR5YyBN8vd5mHoL0+qpA1E8j+YlAYt8Kmi6iwRyE1Qnaw8Gd5aT6E
id1E+VDuusbAtG9EkP5vjFRCtGmS/ZhKocqo/MrhO8UIw5AUrk+YV5Zx4Tyz435vZdUekFQfNlQT
OZiiRdoHrbcLHfF6XKhRoLEHwAPPtnkbHtDf9JSl3hkrspO3b1+5tMTsOwctcJjtYDiweUSzHACb
J6gcb+qphqqdg7G0k3OHRrneNsWhOq8FBZcafA8L8e6SOGSKNrCiByCRSDeMCmPdmCajt3IWKsmh
JG5Sg5E4Fv9y8IWuHO+0VEYC+I4udAm4W8vHTUIp9d8qmYv9qujRRiyNw7Nu8APe3YoxyE6bk2hM
l11Z/C8UfQM0BKvsAUVK
`protect end_protected
