��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR���[{�T���CK��TC,���:�
&��d!��]9�'D`�"9 S%�aQ�`!�6������V�W�l�a锦E(�\gC�slu�4U5=1�N�m��l�9ў��P���B�@+yg��=�}|֦���ָJD�R�x	;�:�E{�t���D���K׏yI�(��"`o�SQ+9�{��]R� ���Є-zLe��%��v��3I	�"�T�m���) ,������V`���q�^�g8)�.U�OU�ŀb+}x�h��I�x2�o����&��5ٝ�'h(Ks�� �رXa�SJ�:�X*Ư ]��LL?�X�'Yn����1�|(C���m��kb����q�X��{���ɞ��J.�.`�RE�<�T�񕝽�C4���u  �Y�����!Fњ#�mv����gM~CW=��ȪV�~�M�H�'�qQ66��ڞ���+E�6�}�ڔx�����,�=Jq��=7�
��R� Lu���� �<M�ۑ�⸵��M���8�ځ���@&�������o�h2i�Q�B�g��|�q�Õ�>��Ն��VN���qC@����}��*��=E����V�ʡ�_��	��~-���e_�+����+ͽhc;.e�E��Ϋ�.s�ݖ�X����C���S�����`b>�)��"�P���6��x���/��&��*n-�每�<����c`Xy!��t	f��!���(��O!��h"�-:[�)�hɊ�1E�t���	P#��^1�����p)?�D�I�\C"�Hx]B����M��n�
��Ï��lO��[�'G��]�L� &R���d��ޢ�U.[����e���>�q�Cg�uh��M��5�����Z������l~��D��?�*���]��ߜ`��xO�������^~W@�ũƘ92?W���a���< |�:!���K�����(W�(q��\z�,9>-�+mݪG:Cp���yc�������Zo9Re�Uc]mz���V
o	�1�?��T�"	#�'�9���}Yqb%Y�2'�
�����Β�4��w��U��f1���&�`�))|*7��/��/���}��sWQmO9���b�K8�[S"��?���;�U���d#��w!����o��#�H�����w�^^��c��,�ob�5�L��gr�l}0���;EplU���A��^i��GC)�U�}m����G����I�>e�;��_��4	��7��� Ԯ�\�Yq�펵���igUﶄ.1�T��ފ�wP��n�͈Q�V�.;٫����kCg��;Ė]�T(��U�Q�T�1Syeʧ����پWXڙZG!4|SzX��{I9���~���	(��͉{��A.p�'-���W�A���p���<�Z�ɐ��N+:�FY��"~	<�PF*��Ê��@��&�� ���}�1vڀF}���<r��Iľڿ�IÕ���zM�FL�h�f�a�Fg�*pAo�a@ӱ�z�Y8���������1X���;ͺ�Zϱ;a ��O�46�ƫ�����I:�$��
؆����u�"���	У���E�>R��Fk��0�(v��ѷ��z��1[�g'�&�<�u 6�S�{��H�����pK>K�5���;�n�$�ʬv� �]''5(���l��UɃ�_�6>-	���
�B쁹�-(�:��W�,#ԁwP/Q��J$�E�?������h��d.b�U�O����y"���/mዾ҂�}.\I��k�#-+�����+a7c��xD��8cѻ�%�!�kslu����H�g�7�R�f�A�)Qt�b|Qw4��D[M����,�_�zi~x?���9smpU��1���~2��0c����/���)����"l���{�W "$sk�Lw���K���:��P<ҙ�,��YA�6�S�1����f���hv;K�Q��jg���7�so���O���xt$��B��c(��ej��}ƙ��ͩ����Y��`K�H�������B`��k��^�k�i4!�d�~�r�9�M��"�'�,0�+;$��q���U�eH���L�Ǭxry�>�W��
��r����/���r�ֹa���EM�.�-x��d<;t.�*���_�;���c�y��l�E/	&� LtW��n�0��F���$�L��%���v�EQ������� ���u�@X|�zŽ>�������Щ����m�Η���ۀq`�D�#p��f����9q�5�f��+�
+�Nm��|&�W��L��=�ho�ۖ��c����r"d�:��lc����c)�����M����׌0��%��Jc��T0C�t��Y���_Ӑ"���W��ǚ�m�zU���W��LR=3��ۅ��d[i���T+OX
�a����F�Z*�X�khE�Xg�
�	��0�BW�BS���|�x��&l[wGDl�9��,jAt]�#	��<�"� �Q Z�ٺ4<�Z-��>�[fw���}�=D�xe^�H�e��oZ�U�	�6�"�j��S�6���rԦX� ������4]vX�w	K��ОӠ��c�;4�n(��o�7�T�����^���|�g�o>�9D"e�IB��u�m�te����mEns���3�"�������O�=@1"X�F$Y�4=�8[�Yj{/0��j7�j�,b����!s�J�_N�+-7|v�C 4����5p��h�(	4�>핔ːhD�X�w��{�ǢNK�(�i�-���u�ɸs;����`ʉ��nRR}�S+�� �1�T���W$	QcvZe93wo�ޒN\�m�%�g�&9Dt���'4u��ӌ������&�p�2��B򢚶tiK˱�!�8XZ9ۚB�:�XL���O4v||eO'ָB�Ĵ�����T��eNU���>%Ln���o�d���X -�7>b��eKA�dR[���ܪn�+uST�+D�V7�ȭP�8,�瞪�Ӌd������B��Y��^��(�O�$�����s�ԇ&�*��7o�f��/x�=��BN����zG�JtO�m|��L�5�"|����7�;R�xr&t/YPI��%TL�QF��6�='^��� y0�㐡hz@�s,�Z����Ν�^1��z��������}��HKI��ݷD�'ghn��K��4M��{�N�K�m�C!C��E��i��^m�2\;i8_H9C �9}���b�zM�4\�?V>JI��28��*�N���`�i
W����5ֱsӈݦ&̒�c��VF���f��QFr��Ǔ�-�M���#���x�v�;V�э+�V2h�5�x"jm�@�Qe����ԟ=�@��ʶ��0$zŊR��-�G�:*�:7��鱰b͡���\B��=�	�]9� ����?�6*�t�l�@��5x$F=-F����3�<�J*�ª��>�;���(Q�^D�)��ٲ���Ϧu��b>o�Y&$Xl��2*17���9���0Fp�H��v��"��^\:�҆�P��z��w����B �h� aG��p+�0b�mVCz���8l��&uH�`H���r��k�(�@��O���W�N�Ѩ���$�����^C�I\<�������@��������?V�H|^]��o�r%݊i%�Ԁ(7O��5�\�B�����xw���m�44��L�q�����Ϯ���1N�U���_a� @��f.*����Z���+i!Qו�|��X�~� �v�O�S�T�TR zN6í�IU�N0mAs�S����2�G��I�_F2vG;?�-�@a�8Mp�UQv⣤]F�)�(�?��"�G���\�J�Bp��~f��)�Z���������2�J�6�[�L\ ����ƗT��}{ww�x}f����>�)w�h�1d4��l�[[j�p���P��b�3b���"���f����x�x���Y��G&0�=��,�x�+ا�n�"�Ȏ,���8�Oa��R�S+��2�%��K�]��-IA�d?�L@��_`b�X�;(rݗ���j
�-O%��L�vU��^oң���������g�;B,n(���B9css��n��HI�&֯����`DF�P5��8wz�Į�P����ܮ�K��O=��¯n�k���ם׸��i�n�?�5�M6�L{���d�Ț���^��ݲG�@l[��[~u�P#�T�r.��y�^%e��Ly߉��&#�"	߈��"����Bx��WA5.��t��]ʀ~�Sy,���D���~�U�mt�F�����A������rK���t6H��:'5�F���M���F)l�Ή~ �o��ۦE	�t����q�B�����Z�beW��Ro}A��	)ܧ���hp�f�n6Ŀ[�����y"�Ep(�f��ؖ��t�*��M��Q�����e�?�X*�|�de���mǽ������ٛ0�K@�7��Ds��|z�l��S��,,�4�^���|� +%PMJ�4���k�!�)�D�I<�v?j|�缙��cm5FW�]v ���;�jx�o�u�a"00��ɯS�7�-�h�');.pE�cno3;������9�Ҳ���O�X���-�����]/koQ��=x٫,r;?
����|^~��q;�8>1�+�w�?0�,�(�m������l���-��E�=#;�R���%��wSX�٫b�0$^�ò{��ѿ�轭@�}�>ny�E�e89���6��^`�}[���Yq��8�(�c��c� 7�Su�/�Ü�*��q�M������]D�g��*���Gȡ)�Up�0Ac���l�,���Sɂ�乩\��wp����f��Xi����"��4���B��ĪT�G�Ϣ+��<�7V�90�`�J���2�Nws����i�Ҹr5�W��4+5�<�44�G�N\�x	��nݰ�oh�$�;%IG��yg���nr�"��\n^r����g� �6�D�> co$E�2_�i�ST��C���w�s�m����S�Ej�^��e�m��~�݌��ŁiR�~i��*�~z���-g�q�)��>ȱ�ݝ��N�l���;'ʭd��
����5N�Iu(A`�G�u�7��j�l��,����`0V�X��Q�^N����`��B:~ɦ����0�(���S>B7Y���������ۖҟW�u�wE��`�7F�0�h�P��M�0���,�-4]\ǉ�w�L�P�FV,���0@�l�]�#�j�lJC�Z7�FET�p)����r|��H�%�%db`-�3�iX��F��'��0�_�Io����콎\9��3��m:�4͈����V?N��(B <�A,�&A�1ݚ1�%����Թ\i
��q3XB��]2�ms����@$��{R
��jƌ(u}�����ѓ]���e`���h���y�]+D�4�>@�m*s�=Ni�i�ա�\��aϮИz�&�+��9�b�\��dNO��P��`�U������S�
���Pt�$���/�IӞ�������E���"lw�(	�B��klT���2Y��%MZB�Є$��W����4
�^"��Y���lU���w��8�H�"�Eus��i�E���2�ؖ0J�#�)}�>M� fԵ���z ��������b3On�������_T?z�#de��`���= X���������i��'���ʄ���v: &3
ˏ��e�ֿ:�I�+��Ԫ���WP�d���z�I�^��;)R1)Ͳ7�Z誥�p��d���n�A=���\�(�f�s��]m��7O(����FJ��V,��-���gh����~J;Fkr�m�cgZ@Z��.>��4>�o$��h��_�AZ&ϳ:ǮGݵ���͜��.z�"�|H�*�_��-~"MO�,?�Q3�ύ9��D�?��$[Ȟ��A\&Ǫ��m��F/����y�8�Y��y2�����
�E����k�ǻ�ʷ��ˌtWQ�U�P��r~� @��BBz�~R&hЧg!����v�k�F�c������Ʉ��4w�K"ȕZt j�c`��3*�e#q���0�{D�1���N�3�� ���2s�U�2ٱ��6��ĜK1�x(j��م�E��)P�|�J��f�4�&���i���}BɕB/,����,N0��)�_�-v�9�JE�Ź�}�9��1?/
�Q�E:���o�<�8u��8�����2+X��	
ם��H�Й���\+�IKNE�Cމ#�3������%n��G��kej���T78	��?���'�gK�7@���d��(��!��X��~(y�%�[���T��$d����!H�oyx.��([�С?��>A(�I�f
���
≌�͑s��.X}�i��X=-{���b�-�2�&�R�?���q.6�/��?���UAYĞ���� ^|1�M9�s��-�}�vR���?���6G��֞v���#9��ua�es)�&X�	��d�h�!����=Ҭ�
�Ű�K�؆���{�kWp*�,���A�[��c_J��غ��8��SE�bx_M�u�L7���e2� �Y�K����9};�U28]�ɻ���|�7mD�V���%0��c{�r`�(��6��2�1Zi*��ekÖ�� 1��yF8:�)^��ܓ�昀	��	.	|��G�3��Fi-s@��E ��6`��ѵ��P�������h�z��{v�]�*�A"r�A!�����0
W�r��)�v˛�d��s���,�~Qڬp�#|&	61�z�V�3�ny<�y���(7s-HVK^�8�(~Q���`+�W��Xz����i�*�i�d��1
j� �[�oP�����$	�[2�a`�\�7\�> )�ퟑᅄ����4l���m���2�m2��#���|�{���ď(%%G����X�J��M�N��I��3r?�!�?�gˬeh^Q$���.Wl�������pM&����<�R���KF���r������Jn(�
Aо�XᚥB�cG7��!g������d�\���A�59���I�@�
��@�c�̟;M�g~�U��d��\p��:*G�{��$9@8�/�8���|m�������O��Ԭ�o�ƺ�j\7�����30��O>`�e}�&ǈd?���uUȊ��n��_�j�#eX�k4��0"�Aޔ�t���'�r������kӤ+T$�ƍ�7`o�K�S�r̂eQg#�6����UL� ��k���8����i7���x�~��L��F���΂�'H���_Tά��&����#����ZY����6\1�}
���*�=��
�!V#�%X���P��{t8YW�;��sո�@;��7PY�j��E�SlnAb�a��|��8�����#��O�ߜ�_2N�LS)����~_�`�^�4�ѷ����{،hE4wGkI�T+|e�6{4D�P�7va�q.AX�8+�!���!⽌�{����Qs�'�?�N��C�����$OEO�!���lؕ�b�RH�A⒚ .9bKx�&�p1:q��O�Qkr�4m3(t��j��y&'��%h��� f]�֚Z���p�m�i�iy�.��$���hBJѲ>@��1�ڮU���Ia����d����u�I萨{�>`�1���.���⎨�=��-�h�a>��}���|bD͆� o� �+Nf)��9��!���#����������ssjl�"��
�Z�����zHE�eV>|��n��Q�r]�ŀE�9�^��aF��Ŗ%Q�ǘau&�9f���Vr�Է�� �I�\M�ٰ��c�s��/y܄/f� ���cy�Oma:�r'#�B�g¶�|��vT��dI�����H6�)�i�t�eOi�����Z4q@M�Jg��rMgv*�T�a�K�0��+���,� �-�E���pCMr���/��a5O��$�ܮ*�m���7󣧉$��99��;��x�!��3���D���r���Nb����>^����pc�h�	��D#1cs+y�=>��:?�h�A�=]����}�ܖ�ޟ��(���,�4�$�L
��L�
�Ԟ��i+�Xl�tH���zv������w�ڿ���S��%��*�!:�v�r��S��=G�(���G�9K���������y�
ʙ0��v�E��q��Jo��.ɠ�������~!nexrb�J�T�����	��=�cHX�0�����D�k� *��#_�(����ʞ�2��oHT���`�[,������s��I?�g��x�w[W[8��E��}��Pv?L�����4�cԢL�����k�lok����]{0���$��s�o�6��������O��yr�~�w����c�Sa�b��B����=&%��	�����#4vv-W�1��m�C�VF�����X���]GG���E�$�i-���N�홷]��G��!4|��o<��ѨG�� ��b���Q��u�18q��y�5��C����^@_	�G��5[��.O�y��V����K2\<�njoo�F�O�����#�SO)C����I���]j'5�?�������+OX�m93/�����O��J3*�6��1]�����9�UO�	~u�E�_H�U�ȢaA�; Dw$�f|�Q�\�g�ѭ�a��in�Z�@����q��W篿��] �|ՙ[|��Тh�&�9\��f3z�J>�C��U�!O�F��n2�c���<S��&qQx��$�eF� 3-���Y ���H�� #�3��Q�M�Ff||
�{�
��x�j��.���w}���4���T�GA�ˤ��~ʛX1��ې�_�`�M�$�FVŕ;Zg�ˏ�=��rq�����m�M���o�h���F�3�T�b_c�}�9�v�ҩջ���6Ա�_���R�{T�$��hҶI�WS��7�U�ӟ�ѐ�f�~F�C���dW��+l�Fpg@-�dYL�x�>3LDe}�%0�%�g4�x�1<_�Ŭ͞�*)���Yvs��jN��ت�����얎�~�Q+:���ƅݪ��(g w�uk$~X�(,���b,��tC�k~	�- =#�`X[mM�w��Y.�l׮��������2Y$��u2�"k��ԑ���f�0:|��.{�&��M*��q��h��G�E�t
o�׼4h�HKd]W�¦1M-��}�丒!��c��8b��ko	�^[+���~�0]ya23po�M�5�:vσA�ѐ"�x�&�� ���ΤCfE1���5B�P��]�hu�a�� -ce��Pa<c׊�c���ؿ$4��j� f ��\�E ��̉��9�����݃���;�#�h�&�C0�C�;:_4+�a�qT�[��7�Hg-#e������Y���:��R����N9�V�mC��`v"��M��� ���QN�k���`;߳�4;:��Х���8Ԏ�s�~��^ɋ׍CߒeYn�S����^F^��G����ޘ������P��Y�FR��OB�=Y�dƥ	f��H����kaUl��+Ih�j�n���9�&�/��R�y�Z,�/����7�w��?��]�C�J^��
SL��M	��R��[�#�P ������1�3S��#�Ď�F2G�r�g� �Fx���Z̞C��OX�y>�_~��t{DN8�E��B�%���C9�l�W$#�3�б�ͷ����%���Iq��¡ԍ�G�B����`|�����Uu0�m���c��E��Ma���FSoԚ�w��]5h*É�2p�2��E�"�iM��S���+_B�%�����9�f����T?_��1(i��z �y�����/R@����)���ǁ�u�WUЕ�������흶���`���$^ͧ�����V
1��s�]��QU�4xv��r��$`HE҃�	ee#ߝjS���쥒�ƨ �}ژ��hO��ߠ���S�JxU����\��y�κe TmΡ�� f���@��"���$q�
0���-ze��$ҵ[� ��c}7�Ho~��������\(�MvZRW���@P D���Ӭ��O߮� �H� U��m䱊� �"�f�t?qh�i���ˈ�w�ͯ��}�Ѹ�/�rl������O�nEhlh��1Y�(܇��L'V�v�H�K�K���ck�-%k�~����:F��GX`ǓȮ�.cf��lȑ�`����Wq��f:� #�&ײH �Rd���'��Fh
��]_�� ~%�Z���F]:��S�5Y�g��vl<��c�(��ZP�W�� ��Ϟ������TJ1����Z��l�FUÈ�Ft�~2r� �Q��M�@���������Lf@�.r����i�����+��K�� ������sg��	=C�B�f�f�K�^���k�Bp`�sbB�l�*.��IS���-�vs�U���U|�@;{DT{Fu�u=!�TVxe~�N��}orn����ҏ@Y�;	Nn��w�h0�IH�gQԖo�;��l7oR,K�n 00Wn�!Cǚ�`֗H�3����m����ѫ�R�oY�"�������̾ؼmj>'bG��O��*��!.�ܽƴ���d�����b#�u�ED�Ex�:�9�A�� �}B�ڙ|��Dj&DkY��)�=I��+݄&f���HĐ�r1mi{)�f�����a�]�7cy��gb	�k���c(x(��V�]%�7ȓ����i�-UG-��\	G��&��M�)�W��ks(Z�z핹��K�/�!tuh���m� Õ��/���=Fc%�8�Ӧ��&�T,s�����R&��=����$&��+=��V5D�F��ENإMc+Xż(l}�����a���ua�91�����_���3�]�O�`tr�PՋ�Y�K��ܾ%F����������o�-����W��%L���A��g�~��"\��BU}/~b����9v1���x�\�h�X�։�����ԯ��s��̳�����d?�9��W���lGҎS�@���Kh��6�3�f�zb��G}t��t(�3*>���*Z������Z�ǻG�%�&%hh���dn��˪l��ƛ�AE����