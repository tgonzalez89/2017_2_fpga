��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR���[{�T���CK��TC,���:�
&��d!��]9�'D`�"9 S%�aQ�`!�6������V�W�l�a锦E(�\gC�slu�4U5=1�N�m��l�9ў��P���B�@+yg��=�}|֦���ָJ&���I��@&��+������.�dx�WH�g���E����'��̯�N��_�htM�80fh�zŢ�%@�:+_`�1X®��iGlt.���\1��B�?�+�v;ꟼ���1b�vH��_�	��d��_ Im�-Z�m\
{I�Uǒ��u�]���̍ 0��%����n3�Y4��@���0�6�d�Fq�B����xVo�˃p-l��=����$�.�?�dH�		����
&����.C��fa���'rG�6�}��ag�g��@�kz>&�ɕ���Y�Vu.ӣ;\�;k�4�[=�zρ8N�k�iǛLOi�Pk&U0�u���wֲ8�Oo�+��ؑ��L��f.qMO�&��ӐQ;ˋ����;%�=��B7d<o���2��3��K|N `����>g=%��wo�n/�������Z�w��f���D�c���ٿ�y�i?�����N���?j����y�so���(,��I��9�K	��g��g��w��J���
�V���"�{��pF.��,T�{�=t��-L�. eE|�����K��+�+�q�}�S��^:֛�<~��oY����� d����]Z|�Q�7�&.�͢y���KdARR�;�x3D	�	 �$ ���-������Z�h�o����J��7�T��"�����SQG���e�ؿ�,�b��=�QF@e�6�g�A�yU����� c��&���׆�C�Z���O�|y�a����:�Fu�k���v�?���� ��$�Sx��s�����J֭:hc�*Z�7�����=������I���6X�=����y��#�-�9����_����x�V/G��i�ob@����.uZ[X�� &Rܤ���<iP���~�Sy?�Z~��?�L�uhv1��h����*_���nVk5��q���-�{D���V����L�p��̨6���fi�S�e{���o�vr��sƿ�|(K�3�:�f�oy�������{R_(�n��XAvwm�VT��nV��U��w�Xm� �C^A4����
����f���#���x�E)�VoM@��Ŗ�X���M�` +���+<�k�?�-(^���5��Z
��{�0�4�܂�%C\Pښ}m�"7��r��Z��Xi��#����#&9�d�\ｧZ��E�{��v"��?��`����6�K{K5q%����)�ӊI�g\B�(	,��#�dz�%ޫӆ��ޭ�7�j�P|�A����DθZ���K��%��6��5z��f��i�'ف?�(�^G�) _���� (�ĭW&����&���c�y� �$�e�qչ����m�yV���h_�Xm}�L�"n�?9k�8u��g���ׂ(�=�1�ʔ`��1O"(�����qk8緋���}��Z�G�	�1�kl�>����;��2P����K�b���:t�^�͝n���˟�ۭE�z�tK�r�f���ǒ�Xsr
^1�[�u0|�S~M���0I�2��cH�'����ɷS��Lۺ�cJl3�oK���>�I�~ثC���,w�׾��p���Y���e|�x���|p�)R�e[Z�7�H{����Z8\�#��<f�R������� m#�.��7�0�l��n$��]���(	�BL	�im��]��º���ޏ7����a>}�����&#*�xb��Ⱦru �W��0��d��`��\������Jվ��I�QmV��ix���1�9K�dl�%����j�(�3,���޲���5p��-TH�������R��Đk�oS#5J:sd��s��o��[�"ǃ�*_��
V�4nU���Z��'�ņ�R)HçI������S��6W�&���ߢkIzz:�����1!��s���[Qำ�7�6`��m=�0��N�k���9ۻko")�b){:�zw�rW݀��N�84���^c�c7i�����`�>�Qz	�K���#��M��d#uȼ�(�dFMMT`�iP�j\�(��+��Mi\��K���QM4����,�?J�-���Q�V4�9&���+ {�+u��Cc�tn���AF�=;P��\������B�v���D�~��ɡ��ȣ�K|`? ͩ���I�A�HC��[���-�^�N3�oX/+�����;ڌ�׹3��N6~���a�j����
�X���N7&�xf�ܹ���'P��!�E�x�� ��`(�z�#�[�G�5�u�+�Hl`@s �JY#���k,S�]��h�$[Yin�ʷ(>C";>�3��Tl6�~!�oF}	�?q
���U/��+>�kJ~ʟS�7��W+'�%�,+ᣯE�B��}-)g"��+-�WG�$4n�p�؝k h�jѯ�M7ujj��?|������$D����q���P���)/��kT�_:�K���L��c�:@>P��� �T^X<L�ڛ㴕�y�}0��ٻA���q��Z
�w��13C%�����7T�č(�~�� ��H��eħS�/�G�b�q��Q0�|W���;���gqC��Sn�Q�M����*p	+,��7\�Ǐ�Q����R��-?DҮ�3 �H$C[U1ح������z� ��
s닒C�w�-/[��Ss���9M���йoH�j�Ua+��u�K�#���E?�a�?̛����(Э��i�_E��w���,��@?�8]V�;�Rg��@�����$3~u^�D-�"��߃d8跄V���Sl
�0:�YД�����v#�bN)^N2S�`���!�&.�є����I�Z�v���I�����?�n~�v���:����|Y�s=�I��N���8��+�|�A(�N�Ȅ��ۛU��^�v��z3Ժ?�?]���x������x�X�fv�q?)pܛ�C6�o�J+�d+X8���t��bt̒yrHF�f��}�q�Ľ��}]]"�j�O`�g�M>8n��/Fk7��5��5 �!���� ]���Lvw񕉮��c�&W\�I�q���M�d� x���>���{�;S���Y�CY�,I���c+��:�CK)d��o���R��Tb[�A�c�#.����r;�w���]�;���(ӫ�p�x���� �2�\�����kc�a'3�[?�Ϥ�1_��^�8���H�Ҥ��|��}�E�{��P�L��q�<��������WLؾW�P��G�
ŷS���oL|�۟�u��b�����=<����5��B�*5y����O)�T��1�Q���;B�ZjO������:�?��Ht��9T�.���)�q�u�X�YQ���bLG&E�`��v�2��3!B>[��~?��w"�;n=�x����j�Ҧ�#�����	�!U��Ԡ�������4=UԘW�UDWHv��Yu,R%�)��1s�e��|�)4^��"8>�n�|�S���y�j�$2p���a���~�u֊��y�nP�KN�0
>�%~,�A�o����n��>��i�Z�X�E! ��g9��Y��1��� af� �E.n��I�I-I���H���ʍ6tLF����7���s�5��R�3A�x}QBp�����r����{����o&l�4j�����#Iw[*��p�!U��l�;X��:��G{����Pß�ƶ�9�������1Tm�PwR%��,&�Р�u�MUf�pY�*H���\�zvb�"u�2,mm���d�`X����pHk�2��'N�I���p��|P�ׄ+�6��^\��H�-���gΤ��X^]);�3��L�+@����j�;\��+��Lf�q��B9Rv���_ԛP�*t*��C����#ր�����r�7�-���E�nʫ�~��cABF�Іg�7W�R1w
�#�g6�S[�?���"g��x�����}k��g�WI���5cET�d���D1����|��+&e����J$���S��[֏42���!%Fp���]� �0�} ��������s���g0�)���W��C8���eK�U��e��_K�o����"��)#�F	8���a���W�K���P�y�:Uw��*S?��8�&υ?�������;U�g�Ϩ�B�;�V^C��3ȝ��R�lA��t�����V�T���Qb0����p���UAE;��F�W��Gi��T�K�_Ѡ9�ow/@5ܐ���؜\O���~�A�ٖ��cAێ�@RD�y�~����K��}�Ѿy����8u1�{�A|�^�1F2��' ��tb���h��3$k75�%z�3�rb��F,v�!HB��`9C؁���n��τ�Z���p�\�&�p��"-7U;�#{��t�'�b���9��&��}��V0�o��}{ۇ9������}qO��	��4��u\b��/�/�5�?�¤�\ꯍ 4ť���`z>�p��O���j�/�}w
��;�����1����W�l=��[j���`��.{���}�����u�|p��Do� �&��gJ�y3 �E=3�4ՙ��A(��\���"�% ������p��c:�T�V>u�$�>R(�/9K[/��`�����`9���)�p�`��1�����_4��z<��2!�}�łO��'6��R��ql4�Z��j`��} �3�_c�D4����H2[��̝\��pE'.{�6H���
�݄��������������j��+��g�-���|��t}0��f¯y?9��T���7�$�D��{������c��"-�]&
�@%泍�� ���=2��yܘBO"S���Ll��Cl�0�����1�Z���0�Y	 �1jO��� �냏J:W���L����P9�Wt�<�K��:E���k�T�=�ɵ#1cM��o��#.]Y`���CFwU-�؍"b���nR�]�y��ux����P�D�V=&��{ټ4��8.���F&���B"�}P}B]4��MՆ��8��k���yH-$d�	*�<bxG1Y� idp���Ω�nN��W:�0�܋'�${ɩu$+���_#����h��F��u0�y�� �������0�����̲Ҕ�<Cg���pS襁�F��b=~Ǌ��1$��BN3���v7ߴ�7�v_a���iUk��k?�y�����7-���i�i*o��2^Q���Q��t3�'�\��/o͗�����a��6��;
Z�N���NWl�F]�����Ř��}���p��!C�����kш�i�&	�X�v�_:�s�GQ�#�D=/jY