-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
rX34va0s0bHll/TDIUpxEBfe4LLb1LYgpHFoLZKde7ffRr+gOpWinwjQPIH9yGAJ8eRInHacwaDZ
PDiwGgQMRy/OCXZ33skJ4R40xjdUm8JJqvOqsMXrh4b5zjGe/q5KB9TSbEm/bTy29LD9KUaHQ6bT
O5ot5Z/2bO+erHFLLGo5NIfUoQ/9XoRsx+VScw/VHRurOXN6y13EJqOBlZUZO/nFuaY5z85ew3+T
oWKwkobIoT2cZFhaM/OSVkkFvu8nKpVjNkvF7PS50x/Hc8G1L+VeKJd6nIsgjLh3mPjXYp38iNIR
ucLVYGDeI5+3OT2q+J+RUt1zEwt+tVO0rZjznA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7808)
`protect data_block
Oj1rtf/GeXek5bZTBWGnTBMbtbJwxWSDS/7RbfMfaO76nIibgGmNy3eBq3fqoGl4Do6smloV9vo7
1pktsHArPGkTRPt4f7JGoMPUdcod2VQzT14aXpIhcYLCtpBytBHbUESaZu3BBB6tJ0JPYnvD0I9g
yFVvfcNkPWw3VBH6iHl3Qkrz5pj7zh1Y20cdA29oivPiiaiDb4RhMfSlgdSmDg6ofYk916ejZZcM
JfTAQhC2qXzNd0J+0YXBuRY0la947GD0FJNqcoTX2ljsfmnTljc0mzfBAyr3nUyYji/gXoaFCqXe
P15e/dACOK/L2aKJsp7PJfrEBYWQUOC3x/4ZDYIcfzhaICJ1EGUSvwlR4zKOVXqMxbA5AgvtiA4D
WcYSlaApf26Vwk4iVm5WUcXkNMbKnzNy60UKBNjMpPhVXTVXQOe7zQWbkO4w6avTJKbjUR4G5NSY
8/AsWR2fkhTFTChrX5hk7/AB8J4FvhOKQ8Ns8AkZKk78AWs3D1x2QSAC6h88iVzhTcbQf7qd0PtV
0K5UHtFy/ywPJaK9U+6y0LaJUptsktfxHXrbhZsEy8HrOBpr6bmvytbl5DRHRc9U4i4j+kJeFlyk
+kFWPH0mzCqbQXNRluRMxtj/R/4p3DPVdvUiVzIVldVpTa/Eo/VybgYT1v1cO653BXEwwdz6uhVP
srxxH9bRx+a/LnXqShejh1qrDBmaJIcrVRqI3r46L6kn7dSET0oU51Ml/UCCEGnH/z8+t80OwEuc
PXFJxSrsWYuDVJ0mi8rjpfQNielkbKGGJd8ewvqa/wdM+vouynN2hh9igFpOMTeZKQnJ/OZC9pxv
8MH3Y4xJbO9ELbpmmCucH6NpoHfCR+SdWZqREYMR5vYNDeCu8sjCtxaB1j8RG5ND4jf+rHmY5eag
1SawlzWGNnHymaVr7H1tv/F1xlwDu9w69HkKz8jc92U/eKdc6qNW1tDKTc/j4fbEvMh/lNWUxJYp
Q+2R/OQHso+Ny+JxLz+Sj1QvlFP22WEcp0NTpODj+eYd3ut0Ad+OF/tKtFJInC64gkGAUP/sPSO2
Or+vigfMB5Ghg8243na+I+DWIs44FPZxJbx8YPeTqbN1ym7GRIxgEet+ZmOjS7s3YfB7+U1h5Cet
YH4O1i1Avxtr99bnpzgE8UzUNZFJXcBZ8V7ODI/DMlrlNw+AcEByujBUataEaB+82aQZy2kRXVsb
mY+buQu8DhBLWIvNx+nFIYH/aFDlIQ8psIujS+6aRnnSomE7y4cItkpeYuMrNyJ5fdfyP61fhk9h
Jp0Xobk/UUiIvGVVjE79XokL+M4UrhhTig7yF+W3iKdK2glrV2syw9kmYQ1zPYKyaiZxYWXjr0S8
VwhufxdrHqxfI7aHFa1lL6X6B1XHWec/v/BGNzQYUJi+ZpXNaraz0xp9Ghk0iNbVs8J3Ct1uxicw
WOBMlHj5CZZwbgc8N3q2TEH2xfafbs3dKIRHZx2X09yfC7rQgynd7r+2NFJfyhonY6LvEvhLqDPz
V0XrssYrxqyYsFLieBO8f7i2FiCyu7GjPBS49UUMxpTjVqmP38Ml9++UPb4mKJ7GhoD3+WqTLH5A
q/n7eEEOvJnkKM7TUf67SURSD70uzCnKWCZx8P5wHObhPqXWs9gR8ZX8HqUE9UEQTKcRN4s6xdNG
LSNoHotkxD2KnJc+mdUnlPOcA/zSjIx5rspua9/TNPQfAhsyj536iXirjqJE1R0FD1fvYh9C0/Fi
Ii6N0NjxwtV1lQktvu1J6N7z6lmuzqyq30YNLFx+EDqQhzlxGe4jzHXKtkSR4Cq63Cc5uvI2R7/b
h+VfnNwIIdNW9xCfGQGGd7ftcXAPcTpN1wONYlo59UMz9VwIohe2QuF9FhReVmA6myu7PhLbLUNs
L7gLBxflfq+JKz07tQ3SoQbuuKmH8E0kPMuIyZ4bDQYNDIsQUXE7tVwnqZAKzPLtDO3+3Ez09f/A
8wt/gxvyC0E3984q5pVqfF6e/X7D8uqkEgPP2rCmBHJIGN4ek2DNCm0VneiqF6GoloZK66qChUFu
134FM6m0ncKCOuvCEW0CCy2oH5dttIhoIlsSmq+153VDwadRgtf4bp1fh7xDanEl6AUPbtxj+ooY
1yqX/P5WUIvdr14U5+Ut/uLfj5tSn4lmJbEPzHUMXAKvWB80S6SRyYKxlGzjXtKkQO/3SHMp0m15
XPDrvZyYwcNTu1oY/5idhFz3ecY3zLfJcIhOZhZFeYUWrTAUUoiAWHjrKOBYBcmwaFRa+dSgiIWu
Uvfuglg+DCMmeLcVqHXTsIh4kMqRWOSMnRsm07MZ1fZhJYuC+oUdyVgUJn7N1gAHxT4lf9EUiYfh
9bkLxKGP1+n3tam1EUze4T3GpqlxMU87ayRqOkQBlsU8T9OA7vtQPEUCYMWdx+/QFU9bs39DGUvf
0bgMuS+jwcpKZJjdN0urh+f4thJviiHuY6S9TdCWyLZBlT6D2MyoDv52Ww/bMF8BSoxxhbWYH2jn
/SkEJzviHK5bb3KWLiWhp7n3d7xkQHrhAcFVIdmHiErWAVtMw6xv063URqYX+f6JL1S7FrAY/UlM
7dKgxf1VLXLeY7J0mXYr6ERFSrZTjYbN6T7CJMuctAGvNOCGwXWbdO5vZ7qP2XzF8W9duab8Drmd
/CYvwIQZlwFusSwkLy2Wg3EHD+sby4OxRbTEydBHoMPOufjsr9GvCnK7aie/xlITpgvenJ2QHnhe
mwBrFLGOELyJN9kGkbxr+abn71d7Ac83QPnEVXrbMEsXT/saQkozh9Qq1+O3Xpk59CGg4EPHVbEU
u+Hk3Bgl2XWUBYWjClkfF6gcLPWOkh8ZKJYcpzUmstxjGgb3mVC3PODD4Xzy7BzZnP0MdansPd3X
g6OyRg+DmP99Hd/5GxHZR9Dv8J/geenBw2sjdzHe4r0C1yKB2+Wd7Eek0wsUsPuNBWa0gicuPPXf
N4hLKhDmubCer6OluLF8lZUDaKkWiIpzHYqF5J0agf1PId1ANA3lMrOpvWvGgDqHC4W/1N/NvKWd
iwbAXXYGAHmv0vIO5XsiTnF1EGEonuLQ9K+KsaXjbAqeSnNj93AQ1cmo/bWA7sTbhBDI9WBkvnS8
gODYIgLn+1CxvynWhMdA02hga/Ozeg3V9LptpnEqqsqsrWE78ptsl/rEhlR4rxjWflnffuDrpUbI
hP18x5Cftzxmyu0V3dOfbYzljgB4i0K8PFGGyLr9/Bey2yGxyZdQ3UFSbSwh6YOS/jRslCaSFPfv
EjM/WSVeJj/df274fFxMbIvdGzrwTdzb7qB455pZCB4g3TJgBXtcJrmBi3Fl44E5s/qmV6J40fRn
VQeEZZZDdAYyYZTbhbCocF9rMNaRS+Z9KCIte8ije6akV/FY2Dcjdl+/Ze8x9jK2SU0YWRzEoy0M
uhdwsh4Zi+HaLUji6jOPRIZG2oXOmJNqBAV3SpV8ltavU6WQ/wr224qWxpyCB9rmyDv6jUmNMsnw
wq17BdXOWUYg0sXRmWym12/qU8S0dSmGgXn8gApkPGkMMdPWHsEMjeNqu+4L21KQagBqE1sCDOZk
ZbOnLrgLlf/g/GZm71+at2/+tdONGro084egIyue6ZnboQgz27h6dLWPrN5RFYMxj+OFx+iGViBH
OkWI8CAYMJgSm4wvjOGPPqcMcsVO6aQexC8MCTsEfoE+QPAl123TyBnQUT9GLHXu2SDoNH/o7GM4
92j1EX7uHp/9C0nxFRTun/n3zDjid2G1CaXWLcraBtNJ/4EzxH6f+GEPE8rdSr5Xzinc06VX7v5M
slSvzSvxx/sZZc/mf+aqwJ6HcRkRI1iPdGRep4FMaMxKwlXxYMHaS2KpyLogeX2US+48bfWoyGWV
EJkB5GKsmELWurzHk1DQqql0ptXPSqjKu7SvZBtmp8J0o0gw3K+GyC3JIO/E0IEtSQQh0q3X+jmE
MCug7U+tpXALyLDDklgmCh7IonlrMybezDSQuQ4y/QlO45BHm4jJdc/Mm50PHRnkGjhiak6hmg4a
ay9zWV98vrFBnHPkhcGmWrVF9u5Y/HVQvwuIHPS+aVHHjsxBj5HHc+xzFXtRSN8nNPRjdaMwXgVY
wlPamiDW6gy5UZ0sxxekQyxJqJbX6B5GXBdgAXGvjJMT+Jfq6zLCjPiyRbVkOdODYyJlBrod1YPs
1T7UiXnGkucq9MFs0iNuC+WRtc5OalSE7S/734/8EYaTUhi+rp3BWngEmaPsGNSbSzijjYb/lkSS
Jc+KACUWEMp839Ei96hISqvnBuMx0Bv369FyZ0IyM4kQGqXuxS/I0+OR1SmPY1vEfCEw0Cw8lLhL
4MaGTzwLEkLHQoEbTZ5pVz9hB33P2NEavjzpwaemPw6H9zoFJNqQtoEQqfiHzUeHO092wVv7LoE0
Q5YFMggEdRjdKDiUDErm67mou0lWbCqZSIWMQu/nsZ9HQu+5DC/YiLLKNFInoXXGiZ881u/w6O/2
7CylG1iZPdgZVDwtlG1aA0F0gcwD20aH3WS80BJFk7ASty/poFiU7gJFc4K5kMQGMl4CKZIe/CqU
mZmbWTTydYHnReYPsaXJIH4pw6k3z4cUE2nD9b0v2GfRxirSCZzMB4XMMXUh9YMVG0WxXEEnIp7G
1Yas/0wc8mZu4iAQd2dYv55KCdXJAE/0Bu2lc13V0bJWAYrZ5sgy+0zI4SoBiBDbCYz7mGkdnT+U
vXDT/nce3pyJIfZzUUhdSDSQGyz+90S/XQw2UAiIELondKLf/DnGZmQSdE4VDsRvsrlF9aQXkfrn
l5JXuUfL2tkyvwgziGjIddPRjCdR/OT6Iatf5nwWrreQvUkzLoxPFAgTatonSAFl+kdzpnIt7S55
EBtaX4E8R5cEQnoAwaPTFxP8nQh3+YsufSQVvke0IUXLW05D0qD3QQi7HCXvKRwp/1MohcEwAcif
z9O8yE9TLaCTN0pb+WFkmC8madL5vNrxOlD4CFNigQAIHDWR8sQTRfTgmVeA1ErY45hLrilxtGTn
XP+2gwJCuyZS0MunTJdyzWC561WKD3Voz9s/sJi3kvjYwasywJL5P4u8mh0LD1LlCb4KTsvEP2Zp
4aDChEJMaU1E2HnrDH3ZjV9SxZoKvoRbB+kWSvFGJ93cebCcznrL7DHN3m+sFLWkKC2nSdNzd9/t
1H/L+RHATIUoN5+/WqPyd7yKsOtItfVQdFLL6I/VGNDosc7CcaXFpu+nZLNOjiyLbhLolwmFV89B
M1nT/dg0N7PfR9J94v1DH8vQQStgVp58dWyR4Ei4Tr32mMX9kNzIUJrCgxs/PxGPoxQoZuj/7SDP
1QQriWNC6VKRlwYfPil3FsM4r2fvJCByMs/v3ssA9bWrFmE+1F0CqifB0Em4tSqpuVolfcqqGYLr
Ka6miPv0g6vxEh6fBG0m9NBYIVWzEPGJhCBIuRWVtVS94IM6MF+bOXs92QAtgp/4Vvo3hRNYU42d
+x1Za34go2/KaqO/J/3YVZec/yUZlmAbVmqawCcs5mUx/wpMWr4rBg31OYUa9Un3FYpp2RowbdQr
FZrXeMWqHBmousIprcAE7c5IXgXDvvceBBh2T21bnDn7xqKCtzOdkIkgYbSC4m7zbDU1kth8nAP6
WmRG2CdeL0Ptz868pgG2VOZho3m87N27yh7r3RKKDFyFK6i3DZikR7lOoFP6xN+VRu/NDdQF+jXP
yJL9Hx6vuR76s5Z4YA+g7XosB3o7ec5zJeqIlhpjsZatk8UXT0ruHcHgrvsmGTwm7712kZf4K21C
eGa8R5nae8z0pU0dE7n7faMAtoK6lAnq87w1sZlFwzYRs2yyiXGVI9uRTH5nRvZY2viUtJhAHHYy
hzMm61ARQTF+x3fnbK3WzScZU8mo0kTh730X91xq9LrTeVYWyHpwGRas6HnsT4w+hEwLkBcYCUCT
GWQ+pcD2mnS6Uv+allhAYy1ZmwkllVbalVFitu/w0YbjB91GYKcDhIu/4pTPcqFqlKtiEAc5T00b
h+NR6SVv7IuIwnO0DGWhgdHPa7mLOucOG3sMWBHSGPJauHdsOpmDssbH0xv+oK3/8IygGcanW4Ek
Q+h7r4aWmsP2hL9N3xGY80SlNirFFi+lNlowrg/VuC8DZibwqWHI+d/zWwNFZzOGDOmWb5RspjGB
bpkZ57ZNfpm1WfPjtgE8Msag61zS6RTA3EpVU4fceZVb+wt5YHmaKkciOl5NUwnXly01dFSVDIL1
qS6fh7OtllfyeYKIZdmggpQ1p9xAH4y5bzmTDgBLcANQUSdH/SGDS76Jr8Opfm6lgS+6Q+pw1I9E
RFcSgD5+xD1fO8Pbvwa8wlzmSDCEODSJxbzVsyOg2b3bthYUCj1p8tSjEI/ntprET5ly6p9xopdW
3lfWuYrMBh1p+DPTNmkcT1fqwrsaXIb/J7qwziAOvlnna71AW8MN31kLftOVvk2YIrs+OjLWLjNq
q7fpmvOd+H/baRALGZ9agRH5kpcDa+b8OhjeXfDLwVdw3zf6fRlnJ9chOmwupNuV2i+JRxtUlyMX
1al4BfAk4L5wSFuQpZNZ1Pspv23x4ZBfLjSAO97fDm6SsHZwv6hnljw3dP8alm732hV4j5Ci0AOi
9gQnZ7xS7iUX2MDDQQP0vwOZ1PPQjynLcu8Eno2oodXf968jZskxhn5jaStAhD8n35s6jewbqQzp
Q71JsV5fy/K6hlM1Hw1/cOuuf95WhUVCPgcFrBsKRFnR7yvbaOFLwJDll3tJFuBFAD6JufEWOOZI
HGySLiVTY0HGDc3X+PyQd0osoSBaogaSBWNwbE8NqTqpOp3AhRmJhnaLE63seRkgtX0xGLYb0aX8
Vaj2NCpkPaZpePz8QCNtxRdKm2xnBbSihvO/ycp17Gi71NtcBee2T4EtPJTATLEg0XflfMJ1+IFj
AjufIkHZBv/UeeSDq7j435pyGQ8j4JNzbYM1Oaj9xS7NoIRbduDbDnYF7n8wxPagMsn8smxC67D0
izzmhjwgc3PylfsLVtcXeDO4xfWuUYiOJexxncgn/gSlWfAy7Rz/Z4JzQcxcQusL/Zk9baiKWUfc
RR2jqBzfsCi92EOO8Vpiu0gi/7G4wYrCgxFOfRCB5PW0lx5jh5EHsU1zybacjOhv8K9HhHBXk2CL
JcpozlVbw0pnUChTLoDbmeaxJYMjoxdHE57lxS9EQPvntHXdKv95DLRepJQHUY2Gx+1OGA5kuoe6
2pOyRAV6vJHKEqB7otOJPMZXz6NBZLqgZy4vovhJFITbLWKGl2f2pf2WzhQugKpBrW/ykCXV4XvN
TE38AHi9xCw879llM1XFMqwL9OIW9qevM3hyqVhf9pEfby9of5NOdj4iUUFoeEHmUJqO/nlI8wej
x46Lkt/j1XfLs9wTp04qmLRg+g/OtEL9sPFjicS0IqpY/Z3wVGStF5swIlPKhlkOAAxg9dF3b5UU
uyPE8/Y2zQd5AJsQ1jEyyjQVkjwXkkcc4gnILH+FmHQRy64NQi8TH4Ea82L5s6Imm+gPF9vodU00
Qz5JbHUj2tVJwGIE35AVh1JEKPFe3esCGntVudp8FNctBjg7HX/G6Gykr2Xhn2OCd7emzDFWiah+
//MJ0jaY+LML/X80xbx3BYJojfZtf7BaNY6jkEcR5J07owVyOUqvvOtF3571ZjBcKpOATaoVVMxk
QvzTvwsDitzD5YjVtdYmtny150KpvUfzxfZfNbgG+XK4CmTzibPH+CG9fqCauaoM4vYluNRG8OQp
Wi6pjhcIZWZu8rQI/kXQUb18oSd/0AQPmSUQ5hToa5QwyvFDMF1mxmXH1dfvmRy57bT21DtGgBiA
w2OQBPLd9I53lswlkALcpU2RTQPb582SvtxFR2HhWrYO4lc7wdXBfGjMGKRa2/Ux3EpW1tnrGTOn
sHT3WQMNUHH5dGqxvrfhbrCQRcTKoU80tq2PbVBZ3irb4dZqiKm3AxrCUGhikpniqCG3Ulzf0FWf
AgMynqKpANTf6bAWu09XNaH6ZLh/YSUUhU/4pBRubGbTIb6+gX+lDFTMv6hf4yNSmrXjzGs/vFQJ
vVizVsUBIxtOBTKbt2Rl9g3ZIrX+W0NcyLht+F4JEsihaJpDg9031ycFbYAlytXN4COX0nAwom6o
iI4NLWndQHBmHwMVU4lzSAkUZirkNFrTIX5PxaSmr8NyKU128uYeH1QhiJa40K4Bk5V8XXJ9Kdl2
UbRVYDVozyvaeAhTVMimIe+iSbxovDagkKuWJoOo/Id/3EurSI5U9XQV7nV2MJDW0+L+zCpoEHFL
GIzNXut+PAY26U/LYpXLEeyVO+tJOELE5uJS4rrgFexT5fhbqdb9wOZiNfT4LWPGVZuqJwQtceoj
F+idHmCH/SJ1iPxkyVSLO+V9e1yM2IWyvLDM9u87K5HQkiaFrWbysUyrfCUoX6ZZAnq+3ulQbj7y
skBgD3SWM5cmzMZwZ54TQrRnVQgrPxJJetFoyDYZXLTQ7//6hROpQFKr8jDmZ5vc0gVuolw0YJjV
0KS2qvNVT0czVoQw+AvpbFdMR0To6vdwfnpWV3xNgIwrsQhIUw80L/gthM55+xDiN+zkwXq0B5wC
MesuDMqy2X4hSrtdlcU3QcdM06Bu33wbYnPHCCFK+pF2MF3mYTRYqJMcyHBdenGdzbCLalXsxPI8
KSSFTjQnwwzI1nkrfwZoxwuy1TFMfoXjSgx+ji6bguidCetti/4zQyagBfGJbzxLwhUWH9OaeCG6
O8xQ4Nd+MYjQO3AXplaeKBL5YCqihwp4iOGnKUENOMq2xXCLYJvWTNZPJSAzxu1ADO2ExqOQSTrc
Y2mtyW2vY42oVVEx0Khl2uxdyp7AW8CSDl+dd49jiyFtKhOL+YKHkA9p7WHAIz3dcWFJFi+6Q9/A
a2uHRcL/JsMTqblR6nIGT5adKdao3XPAgok7govq1D0pz4xJaZFfelJG2G9HRLVDdHuiULNlOAiw
kBmHcwZfy4ruXtNvBXB293lIPF0JXZZzhFegHBlYcj9fraP6A6xLD8pRoZHbk230QFIYLjMbWUwq
KbzQCIccDybjMCh5k8dXRZFn7Ad+sWnB2gzIFi0kCfpMlm/2i9+MEFkoAnp3ildKwQCePrrQ7ZI9
Yxp8oc4Hhxj9MN7EGDcXcnAnF6OW5PDr+vcrH2XmA53ajiqF6gIDF/o1mqI5tfAwSaGrTHrDjxlO
DoH5zp7Q9SHXniNT9pUE/o1reyie4Qi3WIIoQnpLz84Z697mgZqt2hN/HOtQMBCA6TQ9USZB+k5B
eWfUcaFUNTDGHwr6jn8L7OE0xAi2/41MfsK52s3oEc71YFqhRiwjt0DQi39ATFST02u/Zce/lWMx
7jaY+MWuU5be2tMWflfwIe3ynHo0MsPNSoyI8lwmtZiJMsAcYliG6+hq2oEpW8GzUOjnJjLkKP2A
RyzNZc+BrS4h2Ejg1oETGEof6aOZkxqFjeUuRAVl+koK89h9ZuIEPG6ZMIMu2zsnlxAVG/fF8nlF
k4Q/D4iwHua3EEOW3jlrLtgsqaZkCs12ZcIcyjo0qQTwn+1g+7WZvQiPhBFHv0p/aRPRmeR8S5L/
gXqdvfs2//TY9y4N+DB2ZgQS1efbsMGX2+pKNhjvmvnJ+xibvLJV2O4hyOLm5Vgtheyu1lZ9AO8N
IEnBBqc+cAOz+RH63T/0c92w7sT+YVNtMlhPOTZJxjAYBm7N3lNPu98GyAF+08Mzagr3toEalVeq
kX479fIDx7yMIQ4gbrkj5slszAB2WtKfGlLuTAWg4RD67LD2IZSPhUDpce1SkPYJcaOi/4ZSo90V
mIlMxGFLp5mXZ67dkY9TOTlMsESkhFoCo/tK0kIiakCyOyXvBVtET9LbWG1JFp1pphd3be4kWgjn
62GfjIdmk159gETpBgFmwH+0wJkjpi2lMfWWwmwsqX/prDSFF6Tffc0SySxrc6KWTHb+ei6c5yfG
JBIsmWQFk2ypK6/gX2dHxMY38IAeg/ajNmScFNawDBrssfLIoV7Raj4qbVy+74ddZFNBapy3R3Z/
UDHMf1kxuFa/uZcOmF0mVkdy5IEC4vEEmVG60nfVH0a/tUc6S/Tn2wC7sjU9m98uPptZDqsFRKWJ
EYPLyBuE8SBCucstWhm0siqhFhMk8BOYiK0UVTgydtMIfjt6J2dj9bCCM0ZAkbTMaijwkHXrWxF4
2osbXxgYaAG4qcnRy210adNraS/aq3STYrdZKm1vX+oIWW7OHsnnQ3pS7ECDRfwWuStYGm+dk7o4
EXAFFAfSPijY55mkSoQaHTR8vf/kZ6dC5ZXAIGxq69y8C1mhlSTDNOqmuvpczA7ithyp43zAl/16
y4SS9xd4PmHFZEl1Y3fQSK3+3Clh+GsWwqT04hnOB2HCewzNGRTh+JtzWKcLGxUNeZgY2yyWgww=
`protect end_protected
