-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
lPW+pgI5qHQYy5HAHs8ZT4kBP+wEEDXB+46NSjB6FEkTF6MDeIC2ncEOv7nGgK9VlN214jCSWy2c
WF6n/t49/vZLHcMrBPAmfFW5LK1ZCwYorGmOIf8VupV4YB7e4h/h/PdAQgxFb2Q6M70fefru3lvQ
AdxbAtWvI/r2GsgFrG1HDhAmtlT9OKqLfV7nY3d34zv/OzCUPONdoJTydKocJUwRrg7MZem+hEPh
XGoV4IY0GzXJRZJH58nUh4YFXOyhmWJTVV1+oeI6al5UD6aZrg/k5oKJ59y49snz5ljwA+f7j/PJ
7t5m/KMPxy66uFaXbzUtMURf0mSl2tVOH+PK4w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 18016)
`protect data_block
/3Yl+SUQMnNe0jPksUQqi9GEdDeM5o7CvoGbFbN/iUcfgkCn3FkkVszEPMRwlw1foEGaoxB0F9Me
kLKtw2wrFGPA/EywVurUwFztGqUBc40Eoigo2xg3hzyzCziBLI0DcTPCUFQBUCctC9xK1YPBkj0m
bUbBhXa3Bg6PAferqfLbkg6UDk52hSbKDjc3NS337KqBSfxtp40gAk38PKES9LdSWm8Sz2I9nwYp
iIKCdDO6bfKD1ynY/FYLAyliBbW13jyhvF2qAq5khE2OPQ9j1j9Ic3Hl4QmBL55grWIgFR2IMB8d
LogjLPysousjeqzKTpe9DQ20XumimT9WYP4pvsIXqVpFYPe/jBKqK13G9/S4QIzFtTLDFC1t/eTE
SzrqQfF0kx67QKyA1c9LoqILV7RodK4gwK7Yc9H8QR2acuSF4zImsNDYLOcKWvmqJi07/s1eW+l4
51TH+3ND1l5FMFP0Fjn+d/McWtUdtLQ7DDEalTX/qSHfiL5pxB7E2OW54UhSrwELpZAP/7rfv6ml
VinkEOkVgC4ksMU2jBaiXIblqgPYN6IaILvVN68mq01eRL4403DLQUPLRoU5vm96OgexQ4GQOLYT
O/UEFFr46lk7DhMZ9Aaba+QL1TfkFkLCqE9UCgVVsjZyq9LzT6rHZtV6G4FOwbK5NoqM4MNDimdu
JJfY62OAgfxtMJ5IDubywA2UJ8l1STyb+P7IYsXiY2hMAEKlZysUU1Lmu8E8iHo19QzZuBDX5uod
S17kqjR55UzBD5hdm8edSS1HB1gIbMP+S2vkuglDlj26NatBajVon1mEuc9QfLHldOvA9gmGClA3
OwVKFfFB5cLZjmOhH5+PqIH4pkAmCj5zsUY3mfc0i7Ulo2AsnbjSqTT9VfYAJ68OxM+OgB08T9jd
dhZCgbJFStdpAbblRBligjod2E159DHDZXfDHFWN4UME1v/z9KY+4oyEd+ItEiUeIGpMMryu3FGR
mEFBBTiHXtNPfc+Ml+qVUzwT6Ck+PiFEPLIcRgX2HbX1rnJ+349pVYPZg3vC/um480HUNzOpDWnI
7dEhCdmfeEsywtnJo/rQgfa/B0wUK9dft/mA34ZSXLUc9uMe2JElDfWSnXCkuSvUUInyszxT1t9N
DQI9CN8cTSkZQDodyH/YQaH84YjozTBGyWJdGU3QROSMY++wHEzo6Rb3N/MU+zBQpSJle/J8SdTF
hgGSZVokPgfnnRfif1PP6uOQI8mI5YK/TCkJB7JnQZD9fOaYDbdG0zZQLk6sg/4/OmltNIyvRmPe
atMRD4l3st6Yds1aQ5QDZU2A+/zpuIWiC+XozrLpjmgH8O5+ZXdSMpKHD2KA4hPm40qlEz3GoU2F
CjlojyzxxW5tuqSd5hta7m+XHl0dyfgtmkYbo+CMZ7qvkSVRQqUf/LU4JEUX8ni0sOH5LUEipJKZ
YebqcjCVWLkczq6HyFYGYhE4Xek706F5ufguR8xVsViyX77C/4xhLnZCAm+1rkvVIRW8l6kXqLws
rB/uCGn0V6G9Y8NsOOOpV+xuRr9HxwxL2cvGvIRiOfWxFImFvnzOLWWux03VaVM7Q11X9DbkuUh+
PTlBX0Pwlu0ib6PCD3izflG1MPXk1o5Vo3trwW+Kgarr8SI3xq2dA3SnKJrnZTElx41hswW6Zauj
IH8ictcLnHRTRFPiUg8kioVyrG49+qUG7GurhC9bqLgw7Vo4T5sh01jaIyHu3CdS7z69qIkFzfMW
MpoaGyAJXqVSAlrL5mXCk+qXzWoS7r9VBYM+pepIemRAcefkB4kDhPvQWFOZt05wGAj2WYiO1cPR
7Dli+WmiSCP19oDStEvDvPkzu2/iOtdw/o6+IapOdry/5i41JQMqudVl0uDnl5hTIVbUXB0zKrHy
gDs0r1aDzbu1jsjCPxHlNRN8kQbIdIYkREGVg0JWtON4Gzr8WDfMwtTbMYVxF0Fsho053MtgtZtS
jSqXacLih6GBoU5LFk/C//90j/fYDYuLu+clpmgJeI2id2T/0OdxFdTVg04JX01ZAN6BHZihW4Wo
JhlmTM/l4cu4cPxsDFBPZC3fTsv7tRHqApTjCuT85d+Q0h3oX0Qibo+FjtBtszuC7j7Qr+pYW6gM
eTYWQ5BhvO/aKvFs4C3VV918lFBIeqMFWBDpiGiZpAflwLjHQF4g6U7fOsJjxUZXdcHgaq2mhP/4
i3Gu0GLxdvbB5SprlCRgkMYTp4hT/tAcfr2Xn+frYGGoNpJU9kIjAR+wMIS9ekkWlmnl39/osxn3
UOX6TPiN1oK3J606mGc7s3SQxMID1HwdDqxhyVlOmjWiRjOdpVEflVPtNm+YwIMuCakzaLriVmMx
4IWT8gT2Hzu/M7dcBnYH45zHLCQTked0cJnQYVNwjb2JAOtvFrAkseDXzCGXdpTk5gmibTrpW/mP
GOq/DR57EEbjBC1dlAAbIjsdWSPZYqr2v0zMG2dhev5kxTu6NOt5oUujnNrNnIXN+4R+wtpKuNRj
O9+5yYWNwTpVxCGYPHA5GZe/s+rjBpVoN8D52+f2JAjlBAgjTo3KkRPRk2sREhVf4x5mVnCkK74C
GLVKqV78fj4HjgAWgx3odAmEfaTqYpB2VqnOPl1+At5Mh/mI8+WngB9gruk9S79Yjgt/u1mDIvZg
zWfuA+FBzb7Czt3hsV94xHOnGvzHYnWd3ZAdzyH/QARu7v0SETn0X+EK6k9kNrDKVOM+ocmSLhAS
JgF+cKi9LjPL11l6rAtbZNcrzrGJuuruay4GxncpGtXsmSJjF6v8xAMDFrEKsWr7yBEEAEQJGZP3
QmvaZNNKFpZfL/AbgjIH0rRuWLPNd8VQis3OSQkd2Ki9NDJleWMrHEmE2bvq3H5xHJEQSJZJT2W3
PHrx+vJkntC0WbCjUUPQqXaGQhfLvZ/Xk4Ze4ko7cESNjI/maaLdorFwUd/7cIkAlNr+3NUvHtZI
Kb3+UsyomT9E+nofEZYW+fe3/QTpddlhYKoca3eUgKJeVCY6nuaaazxdn9ujqDSWRtGKIlWkg9Rn
egDgiz9VfHqzLBUD3fpa6+o6TV6vDHYLRHb84ZF889OkCMN2wBTh5XDaqoSho63rGoVFaRGfabmH
x78WAc93ngMFGMMIzve5nsjzsA4LG+38o9rX0KSj89w7XUky3hqHT0r+XWGCf+Iu6iP69ATd8N6C
hMKs+bEecWKPhG0EbijYVjKmKNJ4A7SqynxJhM6oIR+pDYeBE1azZqVKX80u5jiMnROiLsburAgN
oKB0+KBYq/i7auWb0doxteO69YKXFOLSfE57V8lgVQ0+UTf3tCUoVppoNFSmw8Iiosy1EYAd6RjU
WlWHyQe6vRxAV/j6NJ2SgWcDdDeHCZ/g82BRwCSWZGhPCrCmSSENnbmqtolx88RN6qePA822lmdl
TVD7avLrjsshwJcpvsMMrQW7cocveL8pUiUMINDl6k19QxyXniSALMV1kFvOkhzImaHfHB80b6uO
qtoaPozrQ5xA99iQVPXGE01yOSWl9w10ffKpJ3cDfEY4bzcmK89vtC/P5IFvCFguncmz3GyBlEU9
LRZtA2sbkYqE4ocK7Uc4nQn8jAfk8n4VMYjVnigjf/pno830X7us2Ps/LLxQcULFSfUx14NEECly
I0sm1qsXThGQr8m63kdAmK66HQV2kZsfg30kJBpw7tjXODZj5FZcEMAGLyhyOsQGl2AuVBdveU6n
cVwXyh0XBdHm/UFjj0YdK16gRhvRL2G1291svirDKkc9NwOd4EVjOGtra4pNXuRAzJ27RUSAIQ6A
O17T97oTYjZH0ALG0GSn1rF5KW53H3FRzLhRayXmTAST57OYYMyaaRqrz/mTDy7+/SJtoEP9z4NM
Eu/wCocJcN3l3faPhVH5zvzHPWqkb6IZxwP3nisMIUNrktDQvvMA+uF/OAcCyofIklt2bDAesLnA
G3+vItfOJLKJfZ2qlxPCu4p1MJ5AzXzw5Wv3oDdLRRWrlF5iDKzPbR+ORpLe8oMr8zrDd1u0sCVE
sO+NJbCYQhRCFbNaZyYrF+FERJJGiCiZ+u0Rb5+0isq8bKRL0/qFkUh4ld5j3yF+HB0iRqTFICjW
+1b2bmDLHHKlMDQGYqhA90mHGmN/WstPYERP7czrv872nApTHspG9UsA9rR70mNScnWWHZIiV89i
Q1Q+BCjo4gnLpNbiBlaLPddV0Inay0rdyp+2A7rmgKg1Z3xkKaDI7ATQ3QfHitra1BNqiUvA1HOE
phM2cGp7y8z+7JmGi0pMf8NGvCFWlUFHagfbK+r47LChDtzexqKO4CnkDkZ4T9qDqGkeSOcTYYmR
h6UcswXWmcoNzb4sTMSz2bQer8hhtT87guCrxIr+qydxvBkrAhxxLcCj9K+AEeT+4GI8dxpRE3S4
xQEwsETCrFJVgNlEs6k7/hhZb6AeJrMK4Cslb+E6XLYumUAXqrTzCtsMDZY2zt+4oLIVpI8QI7MN
TS3MDe2dpIedidVFhdOQXF17vUo7+b/KOAZUmF0FBKo8WNMOen0II4F1Y2KfhE13GOSAN92dsKRO
Yn9SWrNc1yHnUw695B3Fb4KxggChUN/t3Od6VyULZUnPomEj5Wjghs3j1NTgVDrXfIcA//s6njNO
fpiuy2aYG4rocM5wgCrCYBbKo0/VecKpaK+kCNr5wvWdT+5Gj14hAI9WDWZPo042TD84if1kmnVB
eatYvvuApI8e5fD4T+mX1/cxboOKCmOeNAJngWxpOKaizborHCl0sRfXfKrKRE5EVUCFcj/x7HRC
cDni8pblckzXJ2NMYrUwjPKpuMkc8EHoMo8OvBvTuYgyjUtZn+425LF+qKC7hWiRC9pLRjo0uCN4
McjMh+6xVppjK7ZN4mL+8OTEzT3jjblRx19W2Z9D/tJJFAuyZPIFYB0Al9Mc3Ip89dYdJvwuvvmY
M2+OylTYefgZjmX44Od5Lrkovz7LIcp0BgAzHYmg9/l2YDW8i8nCytYKWH1O/sm2Nsp4/B1jQbO+
Ba+nEzdYwMi5cQlYovZiUDp9zvgi02Tfv9ZBqJ8AOpjcKH4gckAc9ikIvjjWgJ2fE4SFWZJCU9LN
T3KDYZCI9xdGqkC6Msl0nKodu0Y/l4IuUrfdRInLJbdzRTSUeFu/fCz2F3lMdsjWAcqcym9lyLAY
fYmlivioGEbuX7vXghOBScKpd6FFNzNt2jYYswfH/J1XLxO5iyZRvUmGzZyfOK6ZOn5HN6/8uwwL
TRooP3PBVQuphAeETgAVR20ohGFl9ObZDblvCqbx6XdSwuH/ES6YlyGc61YOONdXt+c1rO14Xwx1
83NDxyTVdG+1pJwgQjlPbiZIsF9/3VcW7qWK+y8eXdGHAiNIApDNlANWDEeM2OWo3TOsAEv/9bOv
b76HuPbJmd6U8p3NJ9w8uoY5btVM3SBeb1sxESmTCD4qrXFZZSYd8AWBXpkKTgSijZ6rK4X8P9Vs
UGuo3FQA8YLrt2g1lhkpCnwzd0r3jB6Na6aMxbUU4B0C15F7WFWegOUlpqgTSzbbucxJQ3qW1Hde
WZNqEkQ8IScMKEfu7AlzA9O/cpXohjB422atDyNvxghj+2cl08S/HeIbY+B98re8hEoP/A5/xIR7
6JlsGnRHhFQ0DROS+yFB8lziSOOjzaTTSJljXSqcQYTaepRmqwohpfVOF1ANGJ8nGpVMeuKJyNZk
OfRfj1aDCWmt2Vz6cQBZftwas9+D/JT3YTO/RubVgjNh2OZYyFudD72ERyNxuPAoGAg1ClGCVAT1
aUq2p1SEXc3DVFKkNSbhLMSNzkE0mb/jK7V44DueDPi/mnGUaI+7YqpQPA/gWW/5MHg0nqy+CLWu
ObQ3dBBwpvcOGFMnCaf5z1xTGEeDeNE0xaRFqA+A1rKquhm4aniRHurE4SYTkNXyBkl3i0cKv4z/
ihsfI/hL12pbA6FGg5gze+rDYT/CbNSt6AO2QcIoXawHtRlgXTxaS4rJobPVv88Ql6FbTDI71b8R
m9or+bgi16u1llNlW93D8jtXyZyyXLIXn/49ty+RK2iIYqiSurv/ZI74rlnoH4gK5MvITIQbcJX4
0DeoY7brVV/xcSHZZT+7h2pviqHwUp+G2z1hxoYDdDnmFD3TOCb7smYHwrz2upGcTPUWprlvXfsl
ND+XHEchnmzumHctnmlpYVNwiGdkGfKLj+TbS/CpuSkBC9f9aF72WwM/ft4Rc5yx1ldyN480L9pa
goho4m6dnUX8uu2Ym5wL/QcbP5N4vnlSaLQzG+D/Hp1IfwqSI9vJ0NvjapHnbYfUy5kH0403v27Z
b/DqlsYNDEb/yTi3b+vF4WsPmJeuFSyA2/yOnzo90r6nEGqZ70a/9mxIWB7zh1XOFZd2OjTcDXT3
mSsojrUGccgL7YYp8+Ds21t1wv9Tthk8qw4T9H2GNrq9z6sBYQ+dA4g5BeSDSBMjDqcCozT5noW2
6ji++MikiBmEInKNt4HZBILzCDPy6fd2ulykJto3XVqRj+6T3QGH0LUHQldf13/nMw2neHaqeT1T
9PkMxAW+0XEL8kXo6zo5/jAhP90trvrMigDhhQdGGl9fiKv0c8VhYJlsk1BTNosDGA9o6gtdyUDM
qG42AjxggniK5Lm8SHQJj15om/sPWY9YIw5dqMmr/yzwTe+jGutXcki5noZThd5OGMQXKsVQZhFK
SjhSntoTDYA+21T2EVj9SPwz5HooBKKwj+d6cFCvT6ySpFQqWS9ay6L9qtcczpn5PaiYwYr5XUi2
u+GR+ru2i5zh7IzIt6GL69g0YjvM3HVSYJ9q36DrNxl6bVnSlo9NvJrPjc59gu7wTJgKuvLcV7vI
tVH8I+fI+Ey1MNOHM/MYHn85vjRGdri8cAeE96Db8p9F0m8n25FKFUAnfztLdt7yPsl8OrQTSbJ/
b45YC2Iv+TEF6ToKC/kxVy1P7clxEPtIqWviICJj2c81dxQngLxrJVnVqC6DAIf8uUMcqxwvyQ1+
iU7SsWPMHQyXKSBOnYSl+Q0Wkb6xL/ncKf9UAQxHrBZMmwPEKt4J5BJ7/YR6i4Eu3Q/6LIivq7BL
Z0GzhjZN5+VV4VL1As25l5AuE2zBhG7lalbMnWG55RWfqxRgLStX8mW3ueXbNe8IXztMj68Bm7wh
tF79BifC+NtAWwm5C7KYjTj8+Q0CJsnRJ9NDj7qWBOsf/20kx9MF+kCHQQ6Tmpj3iNM4PuTvDwch
QKeX8EDTNqh1tzN3WlxN3s/JDAb4kfyI8v5clRxiTFuJJo0oLFfGWO2lakKkZj2MnPkoIF9WSxul
ueZMEDxT2FtChh5gxVD0y9t/GlmGPNhSxLJsFUE/yD69EU0ovUaU6smKJ7jzuiZR3tOneEQRnnL3
k9JVtHpY4FC7CQ6xBzqB8jnuGTOx3JYIwgavnTAAdbkTv9Cm0OrqFKky1afdq06XRXMaGV0K3cgV
d01OQ7wMkjT/AkoyI8CoPtN97DEJFvx684av9z8z4BQxr5D3Z3zApOIpXsuFg3XHRyTg58f2/guX
nnHBiE4R22u4JcWonYWCGrkt/Eh8Em1u9lpgGklxYU/ftImuW9dwPP/hZe8X1jR8a4oripK1t038
Ev1HtL5XX7NXDUEs8458iqubjdRN+GlyQ2UUE4fjlOy9WI7xX+Gd83ixDlig7gtv/HGThvzfSgzw
qoh7hGfMzCL2gYcmUtDpO3kvjDqLWzRtp62UtTLaVMsRQUpxr4EjLzV7z7uqdw9ylsRqgZJqrwES
tQqb0eEdu3+XahLoA2ffAdmrE58qtOXRZBjDhVrnKhSPTpkoUgK9fdGrk9Jr6zmrMpPI947f5o+F
q4BA3Y6AOQnb0EbYK1FzzYhvdlT/f6JJlTFni6YSgUAxhW8Ly6OTITGtO+ieV/LQ75nJv5z7g2Zd
UKiH7BsesZggagRDISLGXpCV01wE73QlaAhF+LX6zWtzeJOvWNmi8pM+gRrx9mAKUqCblLcOyB3f
1An6PvcXlVlzUmIFzqJy7tcqxi8m4uhus5+Q6tUoajhWbg+g3RYyEKS8fhg2fQL1ODgS93VJ6yn3
x+QI7f4le6I9MmrhBwx5roUYoF69+AMPqHoDh9qFX/rY/ddMq7jmgbQ7GErBcxi2HvpyxicLei8P
fhS8bdeBRNrZVlUPw2rkLk+7ZoEptORagxaI52encZV0NGcXwdJj26mNcN0dzXxtZJ7V9fn7SGr3
kaKlFi2ybF3f52HIq1uP4wKbc5BfPTUTgKbe7lp3vNZNwIhbjmYtfJJB8HQ5UxAiDMKxcfc76bhp
6wyzxpPklce6MHTFEgLPuEf0MHatc8HR2DxG9BTF3Zcn/zpFgCpIRjRDlD4R56wp+1qm4p2qgqb5
bNPvboSBx/9sG1kxuh8ZTvivW2Dx/QhMZSitoHWDboB3+okFB9z6qnBfGg4vJIZVxnCH+Gz1o/Li
e/2JGJpJW0MwQ2Q/RfKT0/8bCtuQ8u6TXOG5sqm7Sryq++h3lA1kMYvSLgwy+ht+csRV5/6v7vm6
7qcIS3bdTDxxx/oVRoa52wdZVG2d5oIzpRx7oFJO7VDrgjKwAv1943qlgPW/McR52mqIRtKR8trW
dGbf1GhNlDYPa/co95Q17+ACAlUFtOosn5xOy1rf95SQHBfpl7dos4Tc2IbdThF12CW9L/UdPMZD
SAT6Q5AG2PxVqlkOspzH0yNZsd78ZAWFEZ1XrcfgQGH+fwrhCwLmAxkZaXe5wCs6geleDfTQOMcJ
Bony7+/lozHnpRhuygzOvlF6to9hgeo9JxTUC/z4cN4Rf6vCGX8kTJryn5k/t/nqnZYwMXkPNTzc
VTe7p2aaZD/A+K+hZ+yQPRan81Xu6dmUu+T9KclvCTkhY38nKWSMM7Vkt8H0UbKVLXUSUVekEFzP
LvpfFhDt7U6ZA3UDNu4pb3VDKBcYK8IgBGMN3y0OFA6g7MgaSwynS9V3YIYM3Ka5xPuEd/ls00Ur
urkkkSxQdKdtjwGWA85bmIA8oB/73ttzvbYLLP5fNevWc7LmI53NKi0ubN6ooj7j7en69QSvdDGS
pRTyIWTU4MIBnP1k/fPswiXSmJNU8iIyl16+TPzPYf2NJRIJwOCqrctJdWJIxS8W+DiOQyIBwAW2
7rOJ1vgLk8gN5QItxPJaQw7t5DiYlyp1p4oQs9gWKV3ujrLWPXONKsqg4z4IVDInmIZMzTkrZiA0
K400mn89/S3bf+RFYUIl8BDAWu2uo/HioCoPI84ZDQe41JRuQ3J/hMayM6mz/j9BL6lzGhPpGgMY
J5NT+WdlO1DgUXIDSOOJCE71ObSubr0h6izhExbr6+12Vg6rfDaJuW4kZMD1NqBR2/BmBiCy3jlU
rU9WTfXdJITObRsRw7PbyzdjGdHZ1X3A5Fh71E/HoOkvUZKrxZ0kiwEsFIFpI1MaP/9Oe/sMCNaP
1vWwE8DKHopK8gRMeaQ7ekz+nhvxQQKQez+TIXIfUSi2M6GLDmmfPW/dMQvKGDThVghbKYIq79cd
jt2BeZsMFzq1zoZhqrqVWQ1uTFgr6CDzPK8uPNXdlqaZTClf5ghtYcQFqR15wH4Zab9mb+X4Tw5E
O6eISGr/FOvrGnRfbtCXtkYNykMy/wMXrPg16dNJNPPmW8iGmDedcSZr9ISLXdKUTSRvWiVrZoB/
FDdESwbBZ/C1ae38FrHNDK5RS+FoD4kbw42hKucqDiCAVPF/MIB9C9Otpy8JQ1AJulCvm3LK80w5
hmoN43WxEGGGVwgGuAUglvdj4ISHWzASg8cdk3pdNDnJm6p7+3dxQ3459ddPPEg7r8c402G1gb+q
EwS/+ehR2fUi8mlCt6Q94Wcz7kKGIKJZeDFU0po/XBMNwF7QtdEczdVX0rYi3zTlDj6m/IbsYi5k
fKiVLxJZGYsWMxblKgUj/pqo+LH83xFKYiHNP/qxnHIQyzP+CnhW12V9/U3A9XjboZUlcGu1hp4P
hhXAtu/R5DsIs25xg6i6fyn1goqQZMRnzGk68a4GWXNpxXRszxiBEX3Vzgbk4MM3uguNoFiSGman
Yy6YRMQVzUk1X9zAWNOwfrrySprw7zymMXXfqnbNylnkx/Fq566fG7zDtaKDN/iqtAuRYOVeGbXB
Ho8IcyIshT9PpsK+two7YhWjEt9L7MM4ShYIhWcs2cWzCeSLAnmgvfw0uJZPp9nwJ104ZvMfiFUO
SV5tggQ1e1IQl6VXb11NXt+pPdqqyqc99bsJQbeKhZR9TJDF4IGz7AtoGeNwQC6J6WDsCAzm7Ybw
FSJleeh42pMSMs5xWnfkdFThfyGEt7wIVmSKNa8w+8Wi81qEC4AOAbO/t0tiyAaWALas4Z8lBel8
FL+3yyjZNhWHd6Q2tJkgiE2x3DfjvhiQsWZUw8yeE3LSTnjPKIu52ICAuueTI7K9TwlwfiF+Uui+
bG4YwF9H7lWNWQjhb5yhG4OdX6Wfbr6/TzxVFJ5m0xLj3WURkL27rZdE1HhQZ0Fyj1i7HNnEcy9I
gv3eiRQPNaTf0VQrvh7lkbyjvf23Yv8S8/XvXNf5LVhED4ipVJBQOIdJ5zd9Z4PAQsxqFhLZTQyt
1c8lIaump7oVKqo+4doDUlZThfILP8x2vXSeEPqOp2JUu3GeTi1GTFI1N9nvO3C5vsj9GqZurfMH
MNR37GtiV0i/pgJcbORQdg60vo6rwJJFd9ZtYx3nH2AdK6mJVcSUxAr1F1ET0ikYSnJp2PdOm8qF
yVx9TBTk9mY8sJoZs3kj5mtJzU9GyjWSJurDGa6pvzoDsCVJPEKKEoBxJ31uGO6Nw4muyLXehKxo
KndOamsLNhf2emDzidojjgicNbhnil9Hm2G+xn0YpU8aCAki0EK6j99pSQsBOXwD4XMsdy97TElV
zjg93xBz3Yk74UtuYEd/FmpPLburmjNimM/o78xvtis4Nmq9l1Og1N30sxvSUZIvzgjzHuoB7djx
VVzUDo38b9B9x2sBr84+AMLUwvgTf3WRiPbYyZYfpvbU6qgP9ZcZrgZByt/5ta+fAP9JrplDKiGS
nxfn7kIT5EyEoMufhDK4Dd1Bldwzqcx2WgJHikLIAeYGhmg/dvhyagbBN3eMLpTd0ZbGo4MVgoST
kyFmxIw6hEUV67XJc7pjYZt7ZW4f+xdse7rSp0UMcDhoOYnTE70zR5BcgESJIDNtUq7HZsbuX+Gw
049iXpDvoVa+I9tV1V+yhr4MkR7QHY4aKfXuGIc1941/BuoOwMIHcnmLHH+pt+gKCvsoqo/J9/3k
adRK6TLmB2E7Gg2wXVSgX9VMfBIxTgY4YViwPccxbRABciLABF4fezECjVO/dgUwuSftEQ+abcef
Vib9hRsgE5KdkX62o8H5mGGBXfxzXxn/4RhIEHvr8xSP6Q9lwJ7GbkHzTYNbBnAhCVSbWxrZ77YQ
wTeWYL+jmWwE0UiqQ6O8kMyrHaPZP8P3sDTOwq83EbpAfylMoR03hPkWOnJpJVtmUMd8oFu+lNoP
MNZgkPP5QBZSHbgxUfABAoABU8wsgyPvnZCWQxv4Ye6P3nil3Ch3JxSZoQmqRPW954gJF6W6Y2ow
csl6dtgwUea4yER8qINkKSyy+NTG/drKlpY8aXbTMTIfZnmGyBXA0Encj8LSS5ZvWfkgLQnLuwAc
RmGABLyiFJT5IMHTBwTojliolBrps+IrupHTGxpBSdq3D1AEUdzJ/1g21YP43sTMkRUerGIb6Grh
rJc72alcX6j+QGajvqPwlnzTtRmzazuUgu4Z/qXUyzJ2B/LPY5aDWs/FmKvNmtjtke3cskMfZ42f
D/S+F+utjoUUyPjnD2VbGwreB+8ejm1aB5ABD+RwUrDMq4ShSeVcRBBTSLyS7EuSWgetmcsiUC8z
4UOwqKp/WjaB3+SkYm/Gh2LzQUHq7bWWPqRawn4ltEaHDSMl+5B+KvY8FtcjBMLO5s7319+ZgQVC
KyJ4saONkaWkFcZfiFpn+Ioe53CM01A+GNXF4ghjQnx5o23LY6qpj4apksBphSto4SMpt9Cj/4sX
9DKH8layTZiV4EsX/kUzbh+IEYc578dBaKB7LFYGPBNRkbMjDxiQk4mbYuocQM3Pcv5tm5x4WhF0
NWuRRDSWwaiZL33HXkkEsopC06emM80NRUXsG8QnYReyZT87r2RbQMXoZDDS3SbpYbSZbadNUvbW
c3NAtlPT+92eVS2B0xNuAPIHEYoZL5BMtQBHjFJNN8RrZJXlx4YKsQmTQW6xwxM3bwwbQfgHcW2/
JNdTgSAtwNBlAT53Byj3mrOZp+sI2tq3k5K0EAjRk8qf82Hx1hC0akshv0mZL5Lw3g8bDS/kCNr0
zOfW1yeYXSjtBDNa29KdjLNlivn6ldPpjJLHvdv0okjKBGedIGDqwypfs95bvau8zaWW3VqUe50v
WtZxaQXZuVReac8F2UZrdcxSH+XEt0H/KmCXN5nN+WmOVQ9sFSKyayKrcLwYdDxPl/zi45AMe8g8
UdLAj6lSFA2eHn+Y/ZGQhQ45QTOELaNzqMNRzqUJKtrYeeT9lFpLA47MO8+1FKxKouHo2L9VfQbE
WQ6fUBQOPxsBuEt/vase5A+f7VAQKtwzISvkm4OLUHvh4zBsRcnDtwWz6Zq4DXqm3mx7iBkemTlm
sSxUfW8NcZMqbQytE7pbJ6B2jKKA2CpQHQgxzcSCkOkvCAga+8BIsKquyAP8trHtZhqjaVM6BxD5
NMYBexXv/5FTxb7JKeKSUTxphdHRPR1KzITXKzvj8Dog3pBrSqBm7UyIAoK9aKZe+aALLn9VfhQa
Q8nfq4EnU9WTXBybMR4cnOe1DzWjmMkhc0rv+unMc9F8//d96hvC3fA/S5sU4HfrqBfwvogo+MMZ
a/1uOkY0jPaMJS8jSwjMjV37WxZRopZsfPaD5a8oMJfV46rVWjZarTQRcC3WAjop/p/mGp9pjoEo
iZZQuZioMnP70F0Hr6gnM0D73n6jplytdpsDAlwRtwGG7c5rCow8zu2DBhwV+VKLMayurEmfmDfr
55uDIafXcffwOyHD+Qy67CBcudiGFPnF3Fl42ObA1Wp2hq0DeQUdb7DuI3bYZ/YQ5XREON1N6j7r
pboK1AUmQ1X19z8G3CT5hSVifI7NBqmHL8h7Bpb7nGFHVJKAa74qjTsHRHbWUae7usjXFr3bbPOS
3iXzlKVFbGMV+/4Zg1G6qHYliqp5ZebTucGTnQnVhgklurcbVYkUMkb5M7mMPVA7hB73bG6B22PB
ImHfEvJdAWthAkIbLqRcDvrU4YxHhe/uMR+kNRMJZ3zIbwLv1kVMj9Ys5Tznno4zq0Qx3klcdSP2
PrR4Z/qEJLSX2axxLHbV8wrOMakSHpzrAEb0MObj5fIcVwBxGJSLmLmXrSzCYJS3dmtKyDdepiIr
h9BhnDzI65q8i34KrFyCjMQxuHMYzn4KYa44IpVnnpQ78jaTYKbvtCiR7diQD2/LZ7nEnaTbZqV1
cXniVhPmnp36n0LXkUHOIEO1Bxod0rZ8ey5+6NrS367oDiLqHNkkWiv5npqucgIueupMs8XjaJP9
JWpwXisUGRFMuAPJDp3x++8ePZXQ2XXFBCSBmCrfVsVvCZdiKKq3H6iMVZTbPR24FwFTxffwh0i/
aPmM2qo0G43quAZAv2Nb86NXipYuEwYD4rZlUQdiAfqabezLQMaAli10r8/85w+/x4dZtJmi0LZi
Ek5TPCsfWa6nWTLd6rq0Vk4LClj/zQsswpMHcZW7AVOONqRt92gZvPhapJSB8jqF7uuSHtFyAf+v
9/9drhx59KNSjcM59Dlz4cR/EjNsw+ZAjGuY7Kqr8evhtlc0E17nSOHuglZwNxErznS9yiiQbJ4q
BRz1hS9irVU3R1un6GWd8yvax4UY0L7H/hdfLuA7ng7FKWJTc1jeNIgyiOX+DDnzqDSLQecvKTei
YhjSFwIlyxE15dYwiZQ4sODvUjOxRH5jPZMTsUFrLjEkNNGXwCAJYxXWpndAbivWo7S+ijsGeoDF
PylnQED3HKAi43Fm1xgWUzBSPuve5YqJw9ZKveTxQ85lQ+8Qr3i8nVRyHTQUfzbMJup9Wrkn5r8Y
HmR8qbq/WWjbI3omtE1NLAiSeMioIT/6FJKQfFxlb2GY6EkNHbf06ByG7l3+v6j30Z3w7iFKUBhz
jisBK5icbRU++ELAjCIWdTbe8Yj5uBBO76f9BO1DIsq2RjKhsNhzW8viuMS32aBseh3veeR5WiX5
iJ4ncZu4iEW9h1EFmsbrPCprbTqAf6qxvk6QXa3hHEp0JFzrchslt+yJjz2FmcUiLDAN1zebjurM
5pbQclNGf8UstLBXlQOp/FvjrrRU3wyOEWp5pkrgvjSkgW0AMKj8kXeOMrP5e5m9EC6r/rkoRxtP
N/6wPlB9psftHF/WIJkY3ejBgwDZJnMk80y6oOM+LvUER7tLO/C3UCH9l5gK45oe42LE9m3lQB3i
6bYv0zvAAfqrUFtbD4IUaKLr+gcNT1UnYd2LArDq8avlwfMwt/k3NC82dsrO8fDwUCD4SD/ADdzq
Mht8qqmakzMnKe0iGZ8u/Hk3gx61O8sGF/scxZxPwtfwV78qrLFVA2QNV3I+PUj55vYsYJ6QN7PA
Z8UtWpfN7tfn/NzI8LVdc/7aAyg0CAn5T6SQTL9Gl0ZMFE5DVvtXspu59YoWrAJwxU74beIyriDf
JICyVu6Gn2c9D7lAWQBCbwMSveNxahbL45j+uxirZtNhsnEJ0uwbxMErjEEULtzzAiDZPQKK9WhB
/MTf9/uUkED3AYr9dQS66S6xQzSssg1twrtl1Oi2+lKOgYkLEiyFCdT+hejfnYHNv2AubBRJrg+6
jRf8TLH2MkwZJeabKp3Y1i9zMkcV9WR9eEoLYe6ENMMaFoCPyE4cwz8P3v7w1OWGbtTz7vY/Rhse
urBip8oOPe6H6qzebHumAJ2GFCzZZp/UeNnWd5aqdae/KBZOoCZIRgnkTggohhRJqsZ/K1O8rms6
6TSF1aGjtKuPhFosR7toE15+aMOfCGShu0feOJIL3OPn9XBnLIjjAu7U8/M6OjwBvXp0LS0NwNY6
Kkrczo2sXHpSFudkj4jhA9SxgujZC265f3V3T8E2zmcDOV2Qm8Ga5pzcnbOY3Dk386M4CwnouBE3
rsRaYzJirkSyxqp0zcqKGlMc9K2poLXB9hgdReyxZh2XOt/o/7nl/bueu4ssHYGDJ4L3wtFabwC6
Paua6RYVWDfn0H4ZOgJv38OyhPHCfxU2I8aVpXIPPprl/QQL7ZE8/q8KYDwqsxXBHp09nl/Kgsuf
/SHD4pvaimShsET3WPC1q6l4LjKhQbzQrIpMq/GwbHdQ5ytdbrSd/zcV7MmptpcXctWRcNQ94b7K
Pa+dDIIQ1crEv5JYAqxvfvGMe6umuk4j93EbExMLv/w7fsxojWl2TR4U70kx3GfJmjtKYF9b9qHG
MA3nU5Ysa5wOMn5bcecVhSxsLaIsqh+5L97+67FH/0tkgIg/6Jw8pLW8BnMsygCsvHQocwnz3PCb
HxoUZNxY5en1m3XREdY23EMi6KCk8i0lWNW4gicwkm5yJBxWQSMrQkNyZ44IbGtumlMTPfYmN6q3
DG5hSP3zN6J2ECSzM6Q1qCqjv97osF2hRJdRMuA5Aq1JaVA3sNULG+we09xtA3DIYRUF8X97CShE
xxRwKbFFiQZagX5LyZLc4gjXC1gR15o9aQlLemdYl3T/VaKvWDCw+nnjqr1QKbASFc5s6ynaKh/x
4XWSFKC3HvzVcLQdK05mXI01JdpI5S/8vp3tclBm9bz2dQsoBAVwTAELj6uyQNUP5vFLmn93v461
p4/H9ylJtIK3Dt9bvB24RE18aWTeJvGKLIYR/QF1YtFlr8aZE4dCrvZbBElRoUr73i4dNLDyPYI1
mqUxvNjl4fTHMNxNFtnVSJgsDGUlyD8G4K7vjmshu3Qy1psodFOUU8PDVOv23Z91/hTzlhycL75S
AdFvSIm8RxCg9kruw2+4I6wSBV4RyEAlc4QoAVFq1hJjYylttm2HgfrR1+aFySmMB8TCtqlXPZ0l
2lhQJfIg19C1pXtc2V5nJ9ZIYCzvoub4KYU4mmQTIXy/tjK5N/6BqSsCjWbhq89scQ8gYLtdOWL/
66EFthkTWOihseXJ4ZpMi0md6vOVfiG30hfojTUwA4IkyOfo4uOlpHw6mG6ka+gVpOGp+AAQ6If9
zFEdXcF9lnNLGanDeXgvYkITxs/mjLZKyNRmYwjAn5JlZPN/z7eYD6Rkdo9e+Z1FSkAvdwvFv5Ee
FeYsY2qo/1nj1uRni7/UNkf2YX7tioNzQL3bmwaCr7w8U2zoas5nEGeVGekkzeTTbpBGuMjDieCa
isxGu7K2lojOVJ6vdjxFVYPyZ9eGLDL8JC3nzhWYNLm6EmWK90nY0g5zJMW6YFO8/PHPlilTfyih
iCuQGtHMphUPmbh1rKdlrFHBzz9rXec7+FwKOGVFt4xzFPRd8nKZs1N9yLXXoXi4wL4pKbwuPeoe
vlJp9dgYHuQ6Fnf4rTnX8LkyRayxZo+1ZAAcLOSaarhOsjBSph9au/73EsOKBU0wYLEybUqp9TXU
7iJ69HAS9ooasgP4S5xk1ayOPn0V3iekGMcvANVtbxQWKEva2pAsnutLqZVuOYKOJDMkxUsQ4bG3
rxojUv631a+oYDwymE6kWGB+Uu6xTs5i+RxItu4RQDSPwK25sxcFRn2YmpO13kD0DZHDaibClMHr
JrpRPQGrJSUfQfN/v0zjeZ82SUuJK7vC++YHllrn5rlGTXDpNL+3X4584AXZ7jtG03vtyPVvajls
c8U9juEk99oy5+RokKTkGuq99tucCmDJEhuq9WXW/aP3EP4U1JnqRe0NGUtrGwo+CxZ4VsKTfMfx
ircTPJS0l3EHgaA3LJh9zfbcmcxlqPScJmz8ldFo5polX7T+14cGDwf4DpaZ7hoGQ/DIC+IEnAlX
LfpRzgf+i0c8mCuiuy0k1nBszcDA6YPmIigN2GI90YeJG1RQHXMPLqIPO+o72l2UQJbMvmlxmNwx
x70kJrk7heth8iOKmC106pmsMkk2WvkgQMr5huigL4OJVnkSz2g7JfDh19MHqw8zPl4BQ4PR1FUL
1RiP8+NB0qbSz9OthnEE1KQE98Y2JOkQSICxTR/o9zBIi2D1qw26I2ffiJyD1TdVYLx8Ln8+Wqbb
x4GVKCGBKSQd5K1FO/7pcNPC6OvCRfEVy2gt5gekVM49N64PkRUU/U4Smx8/4aRfnLjjf9LYVbx6
vnuA5owI10aobFcjAOjJXZ8+24+pl2sZMMLMXmMUf7Vo/jbjH4WwJ28W3biKWOlDl33AOj63Acd7
QpwVgCWMY0q7UpsOOHOg9sM8IaHd/ICZ4CJlrVsCROxmYTkUNZumKxp4g+b8y4AhDIVoDGgvtmA2
MMX/Q1iz62ubS8+MHsiDq3M0sn/mSyOKwCeDLWR9R1EP/4xP4Iz1V6iP/Maz59+u5IZ4Xu8+eVwc
yfInf0INGtVytGSYykjchkSQ9tw7N7RKuStwFZCYVSlNT70WSRDv2C6SJ2EWXFOGhCO6Qr15OKgx
qrAm7Q0+3Q6luQAaKp2zaEjczNS+X4V2nZsCNd+0VC/b0HVMNz5DlGaojgFNJ/5/AltrhYadQ+TR
JUFNFGxDXGtZJTH5NOOYs1+YoKTnJR664NBYBB7w8Cza4FYHeKR+TryNVokUMbe2+TscC9oX/FMv
2aMrrb3j2VoVoWqZR6qGEL1ia/Cy9zVZlInTJuhFN2wlJ63NSaxvajR+XsXoT7tasKeaAjNAQJgO
Mkvr513lYH8YLAYb1qyQDyu92F4U/HsTihVtxrT51yiKJ6MHgmUlyZDDoT0MP2Lfei4zoLnQNrhi
N0krgHwdXi0lvimUcOpSLTyA2TdGSiBDXyaILSODOdCoyFiajRa0zW2C/s36Aa2Zft7UyEmbrBiO
tVQDmpVb1QBBaHnLEGfrDsi2Za0LghoWbSRfRlmnSTH3ZxbgFVOIfom358Ibz6da9iFW81Nxdi5T
ticMrM09pcKL8Ox95vEzvqk0PhMuLy9ZAiJfTrTw7DBIxgXL8l+sYJPoxhINWQ78zwakPdur84FV
mm3lh51hUfL3NSBeha76F3M2ZLmNgC60rFF2hWvROfQJPrjsylaSiXMtbVJCTxYc7ZjHjPcu12Ia
R/tGQJVdBWvysqNpY3m9DF8Z8AeApGdUcc6uXV68khfNj7N7WqSz1RtjGXj3dKfJ0TCIdKT4Zuch
8hhCFA1e5AFvqfLSoT5Uela2vEMdIvuh/AB5OJvTg0/uSXXFDeDNbXdLIj8+Xln01743/mT38st1
IEwmHxNYrnL5hP5/zwNd9F/2AjXnHTyxwKmhKiFGF+b/lbhBg0ziMe9qjOPkcPF2g/krq+h4bl7t
ggvCpTk1m3pZPqs+0fms7yZhou//dMXpkHgnkZh6B4+iDO4CeGonEQkv0jo9CrIT4EvNdnVkn83K
HKjC1wl0wpKy0lY7HUmG/soY3HYyUM0hgAWd1XIrgMHnRXoKF4J4GcVl/LqBCh2ZH8yCiGpRbV+u
tQq28SiXc9PPh86I7PDRYtKC+Q+DqeWnkUbtPhUDuqMkpmfULe3j/7wFWzn2vy//5+gP/jK2oA/V
yctMnDUa0Gb79L96d8GAlLjvJdrf+kcZ6vUJg8xwb5AFo9PFu1WcftmHFrFD2ir2nfEsADehN7yw
NhfJHzUoy1THkk2XBL4RR6S/vjy2tCWwkfXuOR2vdASfP6Myv9vHCIwgVyy5j/F54CDse9RkDTqa
kKcOmMr5rSST6OOua21Kz/zRicSnmdW6Vz+DIjiGtvUNUW3IQwb0FRY2UdwGzeiqDJF2YlBOxqj1
STdA1qbSK/yeSu1Hqsgaf+8k3XvfsF639sVbiw67RO20SLcYFFiLKnz03vrnhQZ/9s7R9OhkgIwO
LZ+nF4K+fGgYP3v+IruA2e+7nn9zkWGScpEGbJNtgzUbu+/qv0ZYxxTe593Jbwnj+yxBQWfDxlGa
ZxJ4cxydiAk8Q0EViP+P5r8xLT8pA7jtLLO9x8CvF+j5mPTsmuqwEzqWelDc0to13QJXWPpvZfCJ
as23ofLcsUDhI97cvfeUPiXtGYr6Tz+MQD2KRs125++O4S5z7p73/AdKgwTZavzltChayOYp36T3
GxqE8AN3qnXgEkboc6zPNvFgWz2J4lRlM47gMUD41GMJf9BRmAHZrebAIXSdU4mtRk5Zaa9MJaYj
4HwZkfocyJvhS6OTPOpm8sq3rmh568Nf84idKPX53cWVIQgfITXWhhqVXs22qfOVzIdAlV9VwEwv
v4MceTV5rsuelYSvy7gDMIAq4xcLuV7rYFt/aTZ1cCGdnT14z/ptG9OPi/KpID1HJwEpB80pSx9F
U9IJjEwjU/G+kLSGpkN9ErdEM+nY1ycpI3SOIzk75R7WhHq9/i0rr5hysGv0U2yLG42WaEfsiwoj
t9LquSvgREjO72knofE6gZRami8Ksb96zS6GHH8R1V0ZJ2Dk2IArhu8QReN4Z8FnyrAoRw1NYw52
uDRo3kZntTdQK0P/Q4JHlBeiRqtfqD0DJpSvct7XWSVIVmlqiw2jKbaE1mElA8U8dT+py2/ctErl
56A/padWxRGrafEPW1DGflr2NcROwjRrusKnXzNVa99GmgYUiUs0b2GYJdEvrG15EDXcPo73npES
BJVP+3aBg8F39oSageqUqIJv76g7arx2TGG2KUVr+O+Wt8oy2hV6gdGbR4j1B8XtY41v/N0t/Fbj
jdFt4KtF9kQUnOSnosPr/MTldH42rNQQqjgkOVylLQJphzG1jozjtG4eUELuZV8szDfeSWihpPnu
+TUjLekal+g2L3Nv6WdykT64SryzMiYM0QVu409BD+FzcbHV1ubJ48pKMdVW25eOIOw8SDInVaxe
o8ECauvA6Wls9Pz/I9FlDCnI7KdbdX8GnY0xOVLP8IFGAReClANvXUb7xBMJ/g7uoBcSVE2TX/JB
zIoLqyTwEtJNnoZW0TVYaPouNzTsO1iQD9N0bzW5rI2L5RwxpVxF0GBBmDmHbi7ISt+WFWbu622t
3m6EyoXZ+1gAXoFtXCdHPnkTKZVTEbAfMNQ73Kc+aVtjzKjak/ceLuFMWCDs32cFyztvbQJw0FDu
VHpPATqNHNzT6XunxjZoSKGAN8a+pLz0jpFksPAGnYfDN2hLsI8HHhGId8XcEJXlZcrOCcmyZW6B
PLlKVw2GZ+MZPF9qSDsV35I1iTbzObA6ZRDjqagmxYDyL/ahjg4bNbPBxOtwXdbK/pItIjA7yb8T
Q+l2vBkisbfiR+NsTqFIsGtrbAfBCtdDM5wNR7gzV0dO/cmlXo6f9VDkQZWhzuSiawOQWD8yhlhm
ocCJTzgaSQELFHSGsuf+DCTk6eytQ+KS4F+QApK3w5v2lSXa/RyVy4Iax9TUEhP6lMSluOweW+QO
F83+vEKKwecGdo3K0vmOyEdjx0lt0qM3uFfnjWV2siyhJsWJvMo7Go4gF427y0cbch8f9cDSWxlb
tjjccGtCJfqpxZqR0L+s2wADOtr/xl5z6zPf2/UE2ox8I/6gnmJPASe0PiEHIhw4KGS9g1dmmqCn
IbdL6PUBPx/FRHiv3skb2I/VgYpYbOALY1OtIcdOnvpMh8Qy1edwEZ2pKo/6BUeYzLE0wkmWaBqY
4EgrSwgbBdEAXYScAAK/+0KLM/KtLyZRvq7flp3mSl6gEK1I4vjVTocvOI3RFS22rbjcpkPzTsGi
IYNoCLyoD5kks2xo2gZgdXaAOU9aPtYtMG0w476aE5+Hqy+Ts49ed2/vWMFK/eBj5OSFDSFdZ+Aj
CHfvj2d5KIhrA7M/j/z9oHHTpkWWe3gxGDKFfAkqaHnXHTVejthjF73ZPTWOKJl1ATeeFeyPgHHF
7HM/V12CKC7cx6d2x+jVVOIpHQas92k68884JU3WmPoWsUVr4H/1qy/H3w8x+W85guZXgW1Eu6w2
/gc17lUXZPRycgdgcBusmjSXNXM8pOV1ygTusxNQJDCMwcERsf8Vh2at8fCo4aUzmdb5Jlbdcojo
unuT+BLziCAAnFHUmOoLN4i/Au7Bsi+G9FxqZG4KT/+y4+dzMX2l//h+Vb5w77KPDsafI7v2R9jC
gOmFo1IJWgy3XkCrNC2TVjcvSdY9yz7lFVo5lhMeAgXBHD63UNekUf+RSXBrqG0xgEMkL4OrAHcF
Dlawq456sEBdaEkHrek8skJcrrOPyTJ04epKlqLRkmrHnUproYjXfB/5Mr0Cb4hF9GNJChLOl99t
DmRTxLaJ1UR/WjFt3zz4Rd8e2fEArxJWzd4rM7sqQT1jnDH14tM17R2JZh4H4VyrsDYTWMZ8tFBS
1aTeA579VEGI7QJoTK65FD9cz187pTsjhpFsQMADs4J674fu7rB1+EAOUycZHypZKTQ7kcW8cOzB
/sUagtz3x3jO4YJMF+Rnlem4ypAiVaimIFqGDKzRzGX8aPpv7BT1CixvKn87KjM7Z9rmHbGs276C
Ho5YUUzpGPuPlyr0BA2BaXgZ0I0LRo83RIrI1CnfrAJMfl7njF87MseKo7AA0V9Skvf11bc+KdiY
LA+OBLPrzIiAKMmfYN+ohQbkLZdQhyLTuuf/uXlWhbtw1DH//pIb6hj0gzHL0AwwFUHaEe9J4sh8
Ul855ypqA5S8lIDuYc1c8ePniDyNjr31XrYNl49iRVLW1W9zTVYuV8IbOhXesGpygTOZHFRn0zJz
Z7GKA2GUilNIH4JlLrP2AHFe73WBNbTolniIhoIIe3oZk6huBH/Fb8viK+MPx2shEpkJNFD3YbQs
TCG7sLRXg27711VWH9AOWa00w0iRk3fhITMHY5eUhe8yGPGZ1Y/L2OYd8dzFYrO5MuVEXmHm5t8k
Rv111aTINRYKorJHk6Qrj5U0rKMV5rYi61ZwC/xx7DqHuAyR8chYAiFWjOLcevBwdci2hTHcuncY
rbdVRS5SzrfdKQsj0sp7Pr0seEpAgCjGyKUg8nRdnQtmYkqKDEoxA2w9mk/yXPn797YbwcRC1Wde
MYThJ6AYEHChqr4qC5bEi+PxuKnve5r3ZmDeY2s0eWS4K4PwAGlV9h2A+suKJcbSrLRPm3x3J+yO
dUgHnt9MeLDgi+kocslfWY/H/30MjFWps4e6d/XJ56G+jLsR0J0xWI+l22PP7rc9+jYrOeP/hOZ2
21CV/T5XIB07Zj5rbecAnnuRkfr5U6SDV7cKjThQdae/4jJ/BcmfR6yMEBX4fIUwQyPhsZgSnpNb
YjQq5ZxB15MGI7Y1gfTfyxI/17paelqLIuFxIQZPTTPuiw3F526q/l1lTeGA2pF79BF2qUCP3XXk
ncVdo6C6lMcRQZ/lU2LmHGLvCeRqF77Wpw0Qq7snOktPAOGiMb7l3X7uWnbWmJ+EyY6XdEnlN9mA
cGZjX8wViQ2aL9Ui51wxIJTlTWFM5g+t0qjOm4LKgLOgjTvqySxsn2TkqrXdlZpHxlvihkYcrKj4
5IFH9SJDbQYT0zxVIJjpY4xOwDMRfoPPYyNZUuPk6botVZ+xv+2H1FDHPQXKixVZcjXY6nmID1Lb
iZ8pQwdeZI+QR9EUNnNUDvQnACkp7pWxR2CvPs6i0cQNfvZFwN4ruYTL2FAzS8Rn0T2ey8ZOwpJ9
saETGrlQagqgCKYyK1Zon+02PcUJsw5dF/bdMjgLd72J+7pAl7p4grcaMDJNDf6YuqU8MsBdUVCY
Co5B+Aw16GtooaBidb6tDFiYhGBN3J/lICnXC+TxrR0lEufrL5OSXczFtoOVqsnSmrSCspxspyPm
LdSm5QT9jK7p6F+5EKSdKftQ198GW3yKw3ZVewlralQDA5dWv4gFDj7a0IJzVoqdL7YOIa0ZwX/X
F0Gg2AMD8gy0I/lFtxD9NSKxnes2PZWrbIs+4E3tRbMHZYLZxayjUNmqHSeZB4lc/ija0rlQEogv
iV8Yv8WT5i8YaA3ihYZOllNMCG9ViAjPZXiJJJBceh/sNusFjj6XHnzYe47nwqXptKbsp1hQ5jRJ
6SExD7JchJh0YI0rHFj6Zy/FIhFCQrb53pfbTmq+dSEqm9hVY3SFdUGxY+wY7/OpjgrzJRSJF5mx
TkTJu8Qxb4dXVM+vF2rRtcDyD5dcOocSwcXohuBcFJY2AZjIWKOMn9UmYmaWNweYvJ7PahK5eBdY
B4Azhfgh/CERuUPMSSgL8tOjHhZHeLwSIk1EO41XOlYS4gHfc2oTNnT0GrnK5cap7SV8G4eOYRio
c83IS1Hccx+C+iIqWtY2MhTXIIoH9q0Te55ic4vLilnzhocUFlejIj/+Yoj6WccADHH9oPp8YE+y
3vBmdkzIz8tf7NbQFn9IsVp0OqmgGbejDGmBkBL6WQItC2Hd/LKVGydOwg6BUqQvq8vMXjMVNZ9T
ndxWUEU5WZ1bPAbGwJ530Z5/zEFVa/7aKuXDg8lAxAQpkUR0VN4prbD2RKzKfH6D/vv7xt2ioyBl
f0e0YXILaKdH60vRyAibz7c081nev/vJsck5BHA/vTGN5h4VF11Umm5Bq1Yw5t3vzmkBr9k7bI8q
UYZSSqiUgfs2S7QMyHvPvfjYnJsGIScFRlPYChm08SB55sfdngqIJfXqFYFBNlJhNvpcimzPbYSJ
c2AUZ9n3zRuVOhRIzAkpzpbPAGIslvnROgama8mQsSrNw+y2D5VEY/sr2gFQL7zEWnkMHVp52MPN
SIsCcAw/TWEo/2FLHeT/F7bYkwTCz1Rd349qUg2CiGJGtjpY5Re2x7cSjvRczO5op+oVExjkTxU4
ENoQ/UYzOA2PpkgVli6rOqX6fK9rOFxs/t3ZkIZxJsDYycjG8oHmy/wzIaUu2YsxhFbu/ZEzuDZU
VWgOhrh1gHmuV6rxlWzi2LM3w+ADBoBCj+L8khiH3ZqfJvEgb+AsSh/3H3TEdmmVbzqSGdg741eu
AIN7z0q+EEErSgqOYn2pDkSOrpTaw5EkuaUgkowXNqV8HjjvsXzGUGqLG8AUNviDh2/vZOHVQS0a
qd6x1Q==
`protect end_protected
