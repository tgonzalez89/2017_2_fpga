-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
A/RvrTRZR8x/vDflLjMRugwdybOq7r4JX165CzPNAe1qezCfODSrjPg3nsV6s2vm9EH3WUwGDfCh
C7zORE7+nDAikO+bs5Z7aMCy/54YcxrXBKt5uqtHKvMHYnC2WPwxoQt5ALhZNZmtlDlux+i/+sDo
gXdl1W7Rl2/t2DWFCoBY7hLWq1vAh3eiu8PbNglNF3nUlWD0Q9DUyYeAd6kxIyNerGiteIKClUS8
NEIGTFH12eM0GGt6gVuTRN3eRU8MXB0j/V8nmhKG8EhMAJK1auEQWvwxE6J2PKYET0mWaj2cnYnB
tGZqyTP3FC4NbpU2d3KkGIbXIR08suERF9nryg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 11664)
`protect data_block
X2Y6fpiwdWoJsNO4Fkj++5mlVQeJR3H8YNvqSelP8CVErfiyzbtY0cS3DDFe7/GSUJcyEGoSkVPX
+Xtrp9nnP7kFr3u/KVkXzozdf+vmp6AETA66GrtP0KRaFoxTzhhmMXjw0nlz1Bs4llJbGrd0uuo9
zP0B+W29kDXBz/sSmPBTQpNPOl5XpdFJjT5+qG1tG8cg5g/NRIUISPdwcJpZF9uYH+PY2x9rAONY
gmrEQ7bXdjtFsQeK4PRZQnYnQ3K1GSzvKw3ixSpRZRli/ZuG3/H0L3l7kDO/9EoDpJWR9JQcBlvx
5cjpYMAYDf+9jJlhlja5vZOJbOnDJkkigBtKxUMSLSKeHxCD98S9nJPojnLzbbtDfSTK82AFO0a8
CCVs0W0qpHFKLk2a4anU8XXpWf3khTCaZGc7+dKPhIWD5NP+7oRqjfONblJrVMVj05Su6Mn0y1Iz
NNdW5/IbRQyLoTa5ORd7Slidu4IHD8mLDSZwGnuk5NXKdHUwM4EWeK+MbjOFnZVwYPfx6Vm0vTws
htg9RTlcjOz8RCybugw0GlFBApUC1dWj4jWurXWmhc0QCUUssc5Z4FkpnDdxCQ5zKdpfESN0jjup
YStDr3Y8dOiUWJrT9FwqykcLU2vdwHoi/SNUgTXpcw7MjAmMoJvvrX2N4OR93phXs1Z+x4LHqAJH
I8vGcQ+eG0heBjW2UpO1oJuCOJ/WJhq79Prd+X59R4PvHjyKWF8R10rPeoVRS1Z/IBmgWOdfdq22
zRizPXjGglncBoa3mn9GhJFyIT4/p7imyyg4q/yv6YgbS8fq7Y7SUEQ97JR8o0nn0GMkqbJvswKT
2RkK3w89gBPOG4LaHcXzg7XApP4HOAbb57CPSLW1jBSempcHYnCLOX4qd/zxL76HQFlYRVsaMkjt
aIsmb0wztSP5wu86SfCdbNod3d8a0ezF7Omiua8pcCsEMFT2NHnGPmDo9r5nxdt/ZaWmepIHe+Bh
EVzhBDZUJML4u4ZutoNvkFWf4CEUdFbFQUnwmMYBYwuc4UyHF+avlD5wH7NuTvZ3XOHjx8RQpXRw
JHsTJ4xX6iIVQJQ5dmJL2hxAhQ2SePCvwSiyBWPSIPACxy8dFNweB90a/t2c0W8ikoN5t3FdsD+f
tAgN89Ijk7sO1cP2mc9QT+8yZm8vnosxHbQnsKmTvcBFaFLOnq9F6As9UH9CrW/vVC7fkK4biq10
jHdg5JD5xhJvBjGyvgcURBKjBb8ZTw4RDdw7DEjpxKjGUPYlmHtRNi1lXvAaOq4+eGxG7/P27+LH
TDTATiQ2M89cunbqBOE/Oy4uI9913bUY3u2mLf1R/ojyDYiGQC8bxRIyE43LGjbgwHrtZvcPODE9
2gbMEWY74fJ0Z1T73ie8sxRU/Re2is828tzOgAz5rVCIwTHjBxsbkQSgldeoNw0sGcNxNkCQew7m
S7ILFUXIEPizffqimH1nUAQZvnP7m0Xcs5VGgCzPZSaxcDKr0Q/IuN5Vw95MJpcvuciMCel1Fm/U
dlg/NX4Cw7fUpcS/5dN4fQk7YvCYH8nyUs7GNZMPDUlDovc4/vi3vEi2ls2a1QqnesZDrjWb7v8f
pYt7L2x0BlcizcM8mYWRsrYVCw/qpjeSDdHohLX5n5MBHY7S48tC6CfRuVkvhl9qK1gHzbSILARI
tb/CAejHuKrO6dX6sGIRf1LPiAPj0eeKpLzTwxCdNgvGHa//nyRI2hTBjxCwrvQf8/gtvNfBpW1j
al7TBKLWFIIrInJOmvtZH0HRwlfu/EYbS7JnHv/LzhJNk/V8yu+PJIYhKq18RJKBI2aJjoZyOMV+
J9i3AKb/dzll2quMKC9A+tGS3q/f8GdRt2INqCTXV5r2rMKzO+2q3vhwSSYEJdyUEsWFnXnp3bNo
04o5N82SS5abRvrPeX5pbFvSk7S/WMplh078lSqFXomMa3tP7dU8vH9fUUO+v2axuHuYzBi9AVxu
luxzR0PkuJXJFoJfxFeQ9bHTiSMu2TgUoHLZ6dQBUiTTdJXRyutizek3T9AvXwr0yQ1M7Yuf1rVn
hUnJ6pfKg8QswKKOTlNBfMTqFVlC7vrCARxhg0So0YSc6MnU+Yx5WsRhWngkiJFSI8thiRbHCQAn
/zQF/lMTJQjUB3qzu5yIhx2/8MNDdZcv//xwtbckYAt2MnKpn6rcnL4iZ8bAUUVZVlz+5ZdU9vga
Ng3NuLkzAsnKfFl2GzLfTPjPHsdnQW1KGV64uXZ19ncFdutpeXW2w6G9rLUvjOlI04CTiUGF6/0N
q5FBKrTqCCvjOsGA/wiGg0d0PIbjHFlCT4U2qz5kXaaMAyyGyKVdEFDdMaoNve1umIDk+ICW5D1D
kg3cnCUo+wT1YcmO1zod0SZYxQkBDdFaTSlD22svkVx+lj8jXpMyTB50D98nUdJ9+T2X2nRmy+il
YJILnmgTaP4WMeew3CHYnjH1bhGnxh0pgkVyzK+L0bpNPOFXxgbjzS8CzXqR39zxn5LlxV/hG2VJ
MAvrXGzOFiSnJvzVwXQfs9tvb+JZrZmZ8CS0jFwsW4wQeA2h08qH1zAGA8Ckl+0IRx341TEEFJwc
myra0xi62Xq7uZLsVNiR2w0OQi34w4ZgVzaCQHO9jtTu8gga9BgxJiBJ5krHq9EtlDqCARIif1va
8B7CXkTZz75Xji3kkqII1RAG9Q8yoKNiPXu4fRKWf1NzihB6cUl7s20UUlcE454ZL/Ai1sKkFhGC
+DwocZ4oRkdCAJke+jICfEp5DClr3MLnUtHsvYqNxyapgXbEGigjw8FwtUlwKZcYAwxAtQq/uKr9
9ImZN2NQt1Kn+8LcYnSjy8DX4z45u5F1Erkb4C6SafNix4BeQcskEFv8ZjQxREvdWsH85NIyX0Sa
xT93JcNOOzMSG6k3KQXoRy8+7kCvGCbpPX38qr51NQHKaMLFvA1y3I0P2dKWM4F5/5Ix4qoB9IDF
qLxio5IUrZdKizcvO1HGKg+X4pBkH2LIUuWrZAk++xAHo1J1RLd7IiNwoVZyF5Opx5bAZSupXSsa
ZzCD6PsL5Hs6yxpAPGnTeyLTRjh2yyyiUNV50fPBHSREX4c/REtALmYDJdgRTgbAaV/wp/k+FHvN
JAtJogRgDSiQL7A0OZ2rJYOyrA45L6FOgjO+rI6IECPMVwXZKQCnrC6eWyKeqcWRVqKZF1JhfLOo
HtGj9TfffI39Bu0k9e6q4LJmKxEwSQyH12P96Rf5MqTd2aIZIJzGEggD66eozCbBLfhJXmDaJBp7
ImEyHRHB2EZTka5U19kwiHFTX6XtkZv37vyUoAmrVCTyPN2lqaXqMGtIfNzWfMuxbQfez5GW/BIf
R6sJEYhbsjhcfiQZIC5B9hxfe9wd8u1PHBhtVc5SK4haJDfBxi8wUDzhb9NInb4/XY1rYlUcOoWL
o2pQEXozo5GfuAbNo6PtE79FvzMPZoYM2KxftPmtuXxF4DC32ndMOAFxheKixHAHONeV7oCfn6Lw
VyjvjLqGnkHmg+6FU253w93Vu+ICdb7s3t3O3MTl6N3trfcGKNK/67E4Y7TFG0UHeZDQYLRrHKLW
S6HBkteitKn94XlvF8WEDjA/5XuW5gfTp/5wn4qcowq7OU3/gXAluX6fhs6K3sJ1o3gOZCN/nOfA
Fwcb29FwVk5iC4s1WU8yop6Cyg+VmyBTCvEbatuuy0s51126cqKz0PM+IAxrJfioA2w9guoq5GXT
HUNvhwdjD5j8G29TBPsmK6L/R6RAuwukaGt8jIrCgkeexhiEB8vz/Ksu+uAWc+R/REPgIdsI7iWN
2iNeSaUFW4KpdTOTAQEE4zgO1YJf4YMU8jcaqAxqh2qQ77lnSr2tV4Bpdm1RaNCcdgUxOJ7TWFt+
gsQI1wkovTjZvLuKUmAGFTA4CvEEHqBPLX2gstjk6m248tDeZiNfOHbGYSl7+qKCQ03bJHtt8Hzi
EdDIt3wXPM9Yp2DlY+VY+OgNqj/L9OS0968tVRaO9AtTZ/BuQ2wB0sdJ+JwKMSuFiRDBf+LtKoYl
rXsudA8RI5xupQ7suodM0OYGLjSW1E0+pbT9+OsTvlnHoRXyeOyH6GLQW5XtBGkUh8iRflGm67n2
MnUHhEXs1xwqjQH7RLhYpFy8AtlMswwnw8IkEXvZc1ga0+g7dz46e6tDbeggTJRoSWppEUes0r9n
cyMYCFYgtPsJyXWDxoUCkH0TbJZH1lKCZcAEv8RxCG0ynOiiS2XPp3LYMnI02SqnVEkS5K0mMfke
xzr+5G93jVq7gj2/uUWOHTGGsiGHBK8jAjZLSzJAh3TEdo979NGfBux+0MJzsD8OfdAGe6g40+e5
pvOP8LolY1yXfJP3naU26/ay+kC8v9kL+v5L5mus/Pl0K/NKnJzYTM37qqhDXxRo7/mg2mYVOwvv
FmLhGmGXymLjq/gYzkEzrLfGfYEPXq2ByNMNA4bW6ISBmD/eK27T/Y4xySgo58xUWDSiY1UGaRAS
uc3OhpF5rp+QeeQjxlISVULF+ZTefEMtXwkrJPF9LaFf4Ja2FXGSO9ezJ3gfJX2BH3FbsLaKMT4K
JP4yV6Hr9pvJroAvLUJoQyfxlJgA/vn1t5gl4GrtTWhSagEghTLZTpN/W2lV8p9POlPKwSTPQMTr
cdEPXF+/P+GHW8I9DsNjvHHBPYbCIV+C72Oe2JjJuUQljP9RCgkb7hq/6kYlDeqMGNNpRRYu2Wza
6Ami/PF8MdtA2mhtoXOQ3dlV6roUjXQLkytdataEUFgCvcR1pXk2f2T0Tlq5XLiWWVzP3Sn4gBLP
wJAEh4xhds3BUy8jkb2MewebT92Xbh3Reqo5lJGFWM2ftV6NfHjofaE9lI7f+eLiKpWzljsWL01W
N3Q6l1OyjyHrteuLtNUQ9as+OCf0Ipj1a47MjZ0Pea+KMiNr3EpD96KuzPJVqLXa9cHFQydhG8tR
XYHMU2HdWClw9b223n2U9lzeUm3y4Q0xrEuhgCcdsMEFUbFAd63dmwsiMlR378pMbXIecwi5haEK
+ZchwaPMJ2dU5T0Luh5CJMgxuyotC1etWivyAtVG4aj61ImFTz48vO0sMUfsTW5M4xd7brErI+A+
X6166F3Br7zlYcxssEOol+CdbrouDzh+pw+p/oPtBSv4ECguJl257iq6K3ocsktL0nl4/SsrVT3P
gQo4q4jf1oJKIHCU9f03+K3rq5eM073H6a/uEebdSY2zw/sFII3fXuPkgZMBXgOfMSIkDvqFcBBn
i68PTXcLFu2p5ircUblxyWnFNyV0LAegNbi9KwiRGwBl2Vn5a0Xy8xfysvyTad+3SDisL/qzTGTZ
m8s+K1wGXbVW3lFvcJ0Bk7pCw7FX6d0VlZvaRlVE9iRqFFa9zoOtAF4qSUwH6jlkFhOyyH8BM8c7
Kta2tl7OjnZLLvH94QrRgDUHHfRWdyhGWEz/gE+TWTwwNSRR13xK3VuMzE4B6WD3lYrId0zdV/bP
diqsAAtzMxuGb8EIwqCXsYp11jBs594kX8o6g93e8qRP50V1qhL3zyrez4yMEcaYO3DNuBFzSMpA
/GK/EBkxDdW44dbcFcbzZQpw7Xuca2CSzcW9jeuT5upurI0RI5JbTUH1UTCzDCxpJiCZANmvIkjy
rfe4XQZFsCl2GaTBEF1nngvwINXkZROmC2niFtPP9LbSMoYJ7o7QethuqGJR3984cAZJjPDG3naY
gWvmJ4aCkKMkoJWEQhrMvyUMT8MgL6bgx90/CtJLmEDMB/oOTDk/pWwTv2LV/+yj84mVn4kRysiC
QhGpMTOo+m4cBqLSgIzl5IJN2jmaBptBJDk0HKH9XEJJcJVahN5Dp0dkyWbwMM+qXoBwazxrxt/O
DZA4tymsJ/YDBoTwDDsq3B/uwQfYjUT/MBc7XBrfR/Y17MUwX3FQ36HYDk8FN32CwxoMQCIDuw83
fh3GDECzPGwYMa5zn+KA088YDjY1k6nl+HX5fxWDeKHjqxMdXYuz76yW8SLVV0yXyeaJEyqUEPAI
WklIvhNpuNrw/YdS9PmYza71f5qvSYCSm8sanvQ+SguYry9wHethZWpYY8QU3kyiDUrUB9Mhf3ZO
kVkrc+pwciGGI/saJXKISIXF0OnuH1pS/gH8P0+0BhKC+qpFbIUH0bovkoEN4v2pRA9R7JnWx8ME
dZQTy7YlZYw9AAM8V3bxQeyWpoXefclshMpIsWjo3XX7z1TJCKNmA+aVMrMWWmaxXcNG1MF6SWAl
C/YxJ/tX5oPcU0u79Jj5C/pYOHhXxnUPIK9nZ6picZCrA0IICUcJ1kdTZnMjW/7mRUrYe+Zrs1Ek
0VyMwJwlaxytZk9v6CZST0MQ4eqMzLk3a1XB5WQbQGk7hR6vvTh2RPnYKKb2wADwX7HaWOOpaNsp
CfFzv5nAes+eZ1tXRyqxTUGUA5lAOWVzd2ByMXd8cud8doHCiJDU4css8VtHO2USwMXEiQEt0QBX
dE/Ry/JvZ7ZDrrsghCEllYLZTSMyFrwrF010LaAaXIYxMDBei6HGX3nZ+05yMoenMZHhxgmknRcU
18Rz6Q7CoVQLIM7XOsdzTJDA31K2DyjzasXiNpo6SXRSl147TUT50rRsJF1I3GQ3x0XOPaS9mn26
aVNGj35fkdM+z5EpjhsZ8py0oAQxYhVRkYVxebVFIrRwBXjAUQVUOt6DYD7KBB9m9DrbJEp+SJvy
IaluZIqcHz2HOC3Or8+CksViJduf47dtwcaPlmNOezd0cLrrMPPDvC2HEZsGp1atey/HQ1nzHNh/
HjRlzbC/m/MEiNp5Gy6XfKUu8bYl7Neky+Mhyr+FKPROJ0fdWBEeMgzSORZo25pxjgl9QxnFCJ00
jrwz0uSPE4XZJBVQXw48DFDQWnZ2bfU/2muA9YmBSCrSx5+MHveO/Hr9umXkMcLqwZXZ2zIefPRs
T2eHC9C/ILAW2z4W5MMQ480W/FJpKll2O07thiEV1jqBI67SCzA0Eu454h3vVKEThTFTk8jIr9xc
IG+awe+eFKDgGEM5aF869k4F4SMAGRlIteu87PyyVzzWfV85dimjFJNOVi+x/u9YOGq0xD5qWxum
jzWJn6p9qMGkBQ7bY0eB1wK60vrB9vNjheQBrXJCVZSFynJkg9SMO0Xx+XuVWHLE1KukHVz02ePS
KFHoe0Pcsusnq4QfxR5C4fkcFx1NaBz0+nL78emlKTsIwqbar4R4SOGPMbQnAk7Op3HMXP9oo5aZ
z2/Pjj7Ou4o541jyILOoMUuXgv1zSJiBTbpAbtltlmwOPrQ+RMe5bCm7GFhGgcEbMxlRDREoGPCP
JSFP3FlVPtHgOmFyjvJvs3++zLCrwu/eP4xWECy+kSISskJWquEImV3cElYs9WZZqZGba1LatAJa
BlSdlpmHscQiWO4EkYpWtDK8/kghcoLYSy4TIpLu/Hr/+4EJ3J/ezH6XX+HS9gk/9sArnKzoEr3T
//ygHqJ4tN1ENUcNABsQxB9wZIYxkrSXPYeT+SvEb9id4LRCn0k50El9VubIFEtvuCDmUUAQ2k0W
u6eVR9O273F2tX7E6LMXBKNISSOIbvaiqA/wDDWkS/vVNUSNqw1xXRA3L4GxDzEWSgdvxiK3LQSY
G459ZEOS4l5VZGackDgr01FY55SUsunKdatl9NGQr65oivgoYvJAg4K3vUNEG9ARL56K1fy8DcK4
HXLP/X1GBbp+6O9qhdb4KIopONjwMVf7l/hEH7u18hZiQjesnSpydCZi/ejAsyS9PF4/4tEqZfig
3bZoSrb4zEDIvLRZsb4QG6WDhTdnsEvP/krH3kor8CFc3fPLcSTyB/kCyEcNMdv1+Vo1f1SanTqO
f2nSqhI85ZCXllxd/YtQ+Ec18seAZ4rj6vGteC0JRqNo+dWngqCsCu5tUKYAjtuFzUPMVViq1nwI
J5AOPuXAFy8KMwcyzpSOON2cKA+/YsWhTAoGZwET9MH8aNuvNSXtllgnH/zVbE65s7gFZ1m8jSo8
0wgTdpLjrZZ6d8KSn44UdWqnuKqViQS8TkEq/U2aAE9JB7YLUaCSzBEn6uVRqKlxP3QTMZelbYGS
qDo+XxbnfVuvJg4FkLm6FDM6xelYuqeUGymlP6tWH1uV6P2hGcdVK43FedNedE91he7/y1uc6AvQ
Pm/bVz9nQCCScvylRo79LkoB/25YuiOwa9NvaBsBQP2H/m3w6oREOzgiJQo97ytIkisPeFVvfqT+
3zccQh0iScKpm2aaWMaJRSlUUL1z6aw1AvcFIq1PDMBXUakrnAHzC9cotgVM7fjvgtX2YCzJgpoI
GFB68APqwYsbNnqozWHuTzJqAd8e8GDclMXmQegox9nsnsNwgtLyEkYD6WTIGTkw+fx8Ngqtw/4f
t0lsT8gdufqKGip6Qo4H0CIoadojNFybfXnoMucPyjwtgbpw7MXvnM22DAwbfOdwWzJxxKa4zmQH
yKE6Evu/h3H8o/wqGdwQhly/uKx+NlYHhKyWB4nHof1ilLW2KPDJjSb1RwbioYWnCFrCQUKxZ3sg
JZT7AkG0aKMXCkTE2Fa3gln8dtYuvTXOMCwTWYlvXlDnDFk1eajUuLlJ/nkpksUUIjFEsve+hIr6
czIvwCII1T9VqdAdipLiWIu6Vx1zLP3cyIhg0BdwbMUx+pZU+jnF74tAizMVQ9cUFtGysagPOHzV
lfNUwBnLro/hI67BtZict/WrwUAE2hkQLcaZQkjdIrNgkKJ+QUpMW2X2nFSh1IsEhXR6C66IWeid
esQ3G6yWYCzhSmCYR5HfkjcJKRTfPoyMjSwK2DwFZxMYmFWzvdQlrumt8R1UYXilxdSDs7EqqZAn
deOPycm0p6xS7eTN1PZwA52ZjgY+GSdUN5q0oTPIp/sUvhVPBkDorWq4KOxsQ6tRv+w4Rrt9yYpd
8g4URLKwjSTC1Xh29BssAm1UUhoDKTrAH+tF/PsJwgbLEkWz01I1WeCE/gfJbl0fBHy/P2n6JKL7
vsYAfnIT2D2nhZLm58/QUpWuQe1v6dezrpV9Fz0J5qUYXz8RZwywqv/P2I+d5TWPzaSCccB5Blvq
7EeZUr67pf3whHi+Kms9MS9khfkB+pzWoF2KUAI/+ckd7j1LfrYYQC2Tp1uFBQRNX1d1La8gEnWt
P1E7lGextFcaLDnN8HMD2okKgCEmpHRfqgQS5FLKrcw8X52sjxLWYCMCS7Fvoz6qAP1JnzfxWC4z
x9XTpmLdBKnkLhqxvqx6yrhxEztZvkK5F0d4N8cb7p6c1WHsVQyAc3tTyZwUJ4g2tR7gWXEiQ1aG
hQG0vN9bDcsysSN1oU/HH5wTk3HWOH8uGsaB0xNMPWN2ghMDT8cJTKk+0owErT4p6tGZD22BuD9p
qEQPktWhze1Dkv9rdwCoAxWbBi+ivNaCqNvRa05gK98eW7UEVc1b2Kx7Gj+7VATnV6OnI5KrstJm
A6NNamjuYbCBJZy+hWPEn/diwsexRV1MaZt5PaB3nMlkx3Qn3RYbemk4Nj2JA23+b/U8GEmGZz8K
l42W7AAigLAs8PDTkFnHLbxnZSymlef1dhZhDR9c0fXO2zt6J6I2h+ie5Q88M7kFEyIbPTBPrmLk
doOcRrJXsyRqeAapFW+bUaJuRSWOJsIf9gYn1+qHbPFI6ebGixjvv8k+uz1y/dOLjrwMp/H9Qs4+
QI7+3Szrdr82nAdEQ1/SCSPRUScHJjaXesHJOlfOsGTl4DZHjooQ79FwIzROskvKbJZ6crvibglN
pgYo9ISSpsGer/bh2Cw1fc6/OLkWUaDCzfhvdxcBeozu32TvQxovFKnvZ9lSYEX7VQB24yWrMqQ6
Xre5sC+HXzUgOeb0drPlNJEfc+CsqXTshvdocU986eeIJkDygym8nXAaVtvMtJGxM/sdJNWnq6rf
HX8aX4W2d7FcwcxQytob8VyVDA6gs/31lw85pcyoxPfoRR3cgf20nxhR0Q6ia23w254oJFp3UmTp
viehlP0W2f6/pOEYfbSDFYZf9s7vk+bTsb3Ed69cohh05HxjCDQVCN9LMraTMKkxxLUw2Xj9f/6O
FyH1+4yby/3ySY2QaVoG0ArlrQJsW7KacatCk49B4R2Iok4HbmsfTJR/N4YAVipsYbZlyqqwx19N
l0l3Dm+lHGhe3el5vU7qQW5qbPceibsNrXAPDAJcZfdS9YTolWVY7oozYnBCxtDtXVpEeofniSK8
fip9aXlbBcbw+0eYdeMhvj0770pItcH8daJl8NitJx4HJ32glPUCNfvy9OzHLNVMXUv1aKY5y9uk
5nazS8ycgMEsmecQxAxp21j1w6RK1BofSDWd5SemlGuWIk7+saVqZwnyz4oqxPnu5ASXe7OHx0SX
WKMrm2l/gM2maR3b3xU3iE0AnpapD4YY0ZIjNWN5qZR0kNzO5KALGIIDdQqhTRcqkkil46V9JonI
jVZczLIeyZR20g7FShU6eiKQ8TvUKzDgo4HOvvS0AtT3/RtuQpc/z7UkrO9cs8HwW4ULgO2r4qsV
xa6rpPF8sxuVPB9nxo6a0cY0QVqJw4ZJeraUoIf5Xo80+mi9u4lbEyWb6noGMmVFj5s3p/sGPkuo
JY+fOrsaEBnLROCBAix4kTGeE2tKJNFUxRL5XqO/aTzjWGt31aIOCxKtWTwFSzLg5Xsm7h+tSjgy
rhh4iF3xdSiwAuNZP//JXP0FHilCfIqc3fTRSOMqqjUZ3F4vAo2C1hCtWG70TzADcXeFBAFrjG2b
aPx1OtT2HFu8CWvrpppC3UJ+6Ub8oiSQnFxb3uCOx8uHdcQcOsYstJA4nbJDSWqJWrTdYTMhE7IP
UYwk9ljWZ6OQy58MtB39aIIE+VUa+TYZ01LF5DMZOcRCjgb+qPSJhOEmVh5Dj6/lb2u8ybyCW9Dw
HZ8g6Gqr9+j8X6DH+lpRxSkYz/EtRuoKRwd3bS2f3+r5wVEfbv2Ls6+5vKkj5UEe9W3FujDQUjbK
kppqDIqsfScpHO7ds07uG24uOEFoCR1T+9bFBn/zAQpobtZiXhxUFSZNGg3PlAivBcR3Oup1e5RZ
IQfbY5dhzcTwtT9IGu7HYKi1PBKL/9PH3PAx1Mo/R446JumGFGwsGYpFaKHT6bv77SZ1X3HIgwy2
0XkXUG20QaDX0cSGdhUkOjZTOmc+/fQ/WVyALvXnG+ZusQ6ZpB3zoyBN+W0d+h9ViMp2ZtzWVpbZ
s7v43DM0yhfMJXcwgDt2t9i+AzpTBtuyF2hTW6F0r49ICnWDc3smwljlyjVr13jdnYEU0Lyw0b5w
KcZoDHQpeX4k1lScrWt/FuWOxOEz3KonQh+K/CpnmBbBPuYktqThgXT/fZPq3nL/Npa1sHYMsYi+
9FSetpX8cSs0zqV++qn09HXiglBb5Csws3DQo+hvcqLrnYcH/qsS8TemHV2Tm7k61QDYKzAf/spB
3IQrlCFtekwk3WOkkEDvPpLP0YsP9r9Dz12c4MMDj0q2JP874lyvJXk0xpV0lOL60TMcZj+xnEXi
mmM1X4eZbhI+fPN09ytjy2xft8+BRSPUgGT4a9mZ8DCT/j3r9+Tk34JlsvOZ2HlJjJ3Y/7Z6H+k9
Rloz9qWNRXDpRTsiuCKSGp0CvpPGNR2gltWtQ1lguFUXvYqcvmq0LddyGjocE6wYtFXJgM6VSQeU
NrnQ7el+zs2OoOCDXOYheT3qIE0en2YibreKOWnaMn141RURSaHTgbJ188y7tjB03EgoS+7YdJVg
TFT0Ar/zHRXWY9cHQgndxHpoErGuPYHP91d7TMn5hhZNKXQ29EGzhnMKJQPavtUeQIZwcQ9KWXjo
pelvdl1lebAafh1DxXTboNfdB85zZonzhdkAwLJi9BYbm8cNmDSrlcT/e1KOjWw1J48VPwxifUwU
KgEfQ4ynNvjWl8EUarVpIroNAEkvHajqMcph3mA3rz47sa6TkL44jAmFRvAgc6/U7O7w3yfwVtvN
0fjwK0UAsjcGgSbic27JGhdsiWiFMxKC4Wa/s5Ue1D3ywFngYNvcNqpg7+ajeEYyCjcGgDVtlP4X
2/nFyDv0jy1Y/4k4Eho8e0Ax97GUrTFmEpsk5Pe4gcsfgznc2omL4oRr4CG+LRKLb0YJg9EvulJO
1bNbxCDc2sP7NX+s7nKr10XR+0xy9saESB/87M2PGXo+N8tQO2n00ugiNzWfxaeAai6KDDi5SXW+
RBOoHif6qTaAguIokvxgXppklUwZR2k3i8Z62zki8Cra4v3/lw5pGvh4J0uA1Nur8J3wJSpzOlVv
uQtnjUAXhYZSl7FXgrCWnGmin7K4aVoDvrnf+VOo+F5aHK1psGLtMaZPz7f+BOg8Jcl0Xh7gBeAs
sCWb88AKNVKrPzfAwscumX5KkLjXnAnGDptU//vatM8xor8yu1Rt2P1ui6x6z6/IQ6jdnxhUBPO7
d6NXxG6ObmGmFOr9HM6FJ46GHFRkHVVYGVzzTrXZeD/leuGa8mFzS6lTlcri1KLkNa37qCZURwTg
MXpwzXjIwmXQd85TOHRHkWVIz2aXRb2QdG5k7tJL9e+E34jiIZTHRTO66Z3AZNrARknjncfMoivb
PTLyM48Mm78Kp1/V78S4gH/iLxFvw8NSRbiiRepf5jw+117RGjCvFu9n8wpNBX5pmF6npmt1V0Eg
/fOoh8+UUb4743Ukf5m5ByILK0fGy2lZPhKV/Hc3xO1PErF+u0Z4fQT9OIJv1SkCqFOGmoVOVYwK
Ns/K+OJMbkLczv/Vnva7t5thPVHfzThisRhbESOioNhTpSEeC9zuhZ858K/rPNq6BX5HN5J++Tcy
ITVsAe1X8t+x3GT6aQ5moQkIbfXVMSyx2zvVPzWBGAV13LkjnTY3kMQ+QQkO5JLm4kKCqeIpZx3f
39yK4zt5O4bId2PHID5aW61jC6UHz7CWZzjzy5MZ2yNgcjxHR6SuLKdZeJ1ixlUTAcvy8Pm3cGvo
530OI/KI3+frooJtPsKpSOuVar46WBjxmo/jrLapbdZYsGu4TJ/n1ZDm0zxyZkAAziHe+oR86uhY
qui+66tt7Dy7XKJR412Lw9b2dmG4+Zyk+LtDLXOAZzRYmU/+L5scCXueRbxRY6h8xuShDcr9lI7W
N+wPYc2YbgTeoamBRki4anbtst0TwyRc9C4dmRh9gPVF6Fk/LJc7ywwLBs5mZonknYC+n5uI2lcs
cf+/gE4LScW8q02OxDKDGGXLAbSZ8IKZdnqxrgtH0muQIlAQA1aw+sxrv7BHtsIwKZiId+yldwkx
xVtT0LUR8DZUa/s2EqhVRnQ9fFtHFhMFFpgNlQ8ipUhy2HKI8etkme0LLRc02I30W0yruBVu95Dk
b5Blf3YxlY4gzr4Tef1GkQfyMYRqjrHBv6cp5NRZpidbBOfz59kDdvt33AsJd0b7kEWArBaPoZav
wp4gLlgjiPnfZ3W8vhfSbEb2K0H2+r+d/jPIvhSpISm2m0mmynxIqGnENvWqVnft7ZMVhSnDSd0N
YP1hQBXk36oL9CBGSce08vNFXGevbkVgJpbR+dzSvHXN+hxKHCTUQnTNcuWDlb1RCVN7QZp9W5ol
Agrpjju/TALA4uqb8hoN3PVAWJ9PI8g5uxYy4aN+I44/hRY2LqnSGwtZhSB4sq+OE5VI8drox0OH
QEt9WB9fSvEOMePuYQVbR1MEddRdc/u/wp7u3knS6ifNDEge0Q0//pbkpSWbHMQuN7a1wInOnuEr
fEer9FKN/z0W2+fprvFbEr1hhHzyI5MHIv/Rq2FGNJX1G9l9xn2MN8iz5m79dD3opDPocfP2jRS6
jt3ZF4yhChOnjjCpQ8Wq3QbMLSyAk/1IRns+Ot0w8fAMNyn96KvahyJREoad+bRWFow7Vz0qooA/
gBWpdByWAHzJwj+6iTHiG7mXkOJLZfHkAYd2FOTlqB4RkBZiM1FSUUptJ8ltgQhaUhpB5A0CQ91v
LCMdWbSI51t2UJldt/rpXGlS1pyEMnpXU0+e0sQwE1S/FtjqBLrb08TwzfEgbsQo54C81grMd1mE
ievZNgeEnhDrnfCbc8u0Hi2GAnX4EVVt8V/h+5dkqJWzL+o0q2/4eGIfVA0he9Yq79d52YchaLb/
1it3h3MIq/qZZgkDSkzfjJiZ4vUkZ5gaXltzQ9HbcCDs9f2a81julswsVPinSjZd6HUXpdPZdlHi
jAUheCfbtTGrE/CAXvtDI+/PsHmRa+WoxmwbTYP8lmqbTetVNNDUURDr+h9QBi9feuK681kKvGb/
CAV7F8SUuOuWP7m+6oAVpZpjNhwAdOHLMsVW5mHM5XrNoQlfK/8c2FScu9sGVxDPjJ9DbzwoOt3z
mBBxU9OQXwxi6GQ5IXjKbKJSlxR+cNj5RUxcGG4e5yrvWay46mkjB+eJWOAtLSaXVVvYEl71AL2L
4tmN56pGE/X4i8gEmppbHd6gn9EciQbTU2A5wJA2wLt/q51OIeGrY3HAobLzCvkTfXaJMiNQ66G9
CKbNR5f3k3Qq1cndH5d0JyzOd3ucIv6geP7E0wqvUfnFv0mVh7yqg75txjTASAR1+xwa4lYL2PZc
33GtH2eZ4izE0kkJ7LZ+7igr4pro1zQ7zQU295LgyNcCeskZi9QrirtqmpkWfeiLHCe0IqIiLrSV
2nmdMkXS4C3/0RMjcWypjSPZt5NavCL250ViqgHdICEFeC5e9Dx37ztcxmoe0g27jlz7bhOy89JJ
YnREJPDQ99EoMc/koDNy9kRH7PvAQKoolOUCdxynLqcc/oXJ4gwcrZUry0Y4immx3G+JopCj76Dl
x9vIIRurpWyWmYt9jLvtj7DJgkAm3XAQh/Ij7NIqq9dhYqKbX322V+34uPJwYsDCGYMP5v9Q6gHS
TnfqVLnb+r1BbygEyYRUVn2RSQNZ4Blm4AnagIztBHC5BTqZCVz5qnHijbX3wqtQeVC1Eo0hjhoK
d/0+CNj7ini+nwdWlpWQBijc+vrwQmQNWx+EAk5fkaKekS/veB5rwEzEo/tc/4D0JyZOhYl0/2zI
nfoII7/Rgba+oEluRzKI024Ruf1NccNs/buQ2j5BoUJEeI9oGXgQy9Ne0UoKr34iuuhfs/T8MGRa
+u2zFHcWXM+HuvJHJo0uMJx889cWYURDoFglpbID8vm8wOehcvEmmRX8Syf3dPbasXj4CHpp95Qp
NhgejtoX9V6LeS5lh5FNTeacb77vaRSn42nYdq6YA028PlTclEDV51QCdx8H77jaGzZlwIxbYpmC
tyVhxTtqg6yoNUx/x0icwlxU3MFBwn0i/wWUoYqghb4FnuHC3dYO+mjUdtLH0jxuCUayqrhatdWp
pBytt2WgRF8Zq1aDVMO4k07mp970war2LvFlZ7Fji1wfGFpzfChBOvI9LSVM2TIAibIrlf7e5Fww
/nkzFxhIZOPiIlw6cYPjGfOBiCMh1Mk8WcIaeb4N4NnLyzPH2HyLzer1EYH28VELq6z0N7RbMX6z
c34UaAGhE29m6cNYNJNSY9ovfASlkddK+iAXYWVC4ChRkwtoWzqAq2lHUt06rOw4iZeHu7VAQnZQ
Brn+4Ax2Asa9v9fJ60V8URJgBSkI8PG0d2BwOT0jWcZFN+DT
`protect end_protected
