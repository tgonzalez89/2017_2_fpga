-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
fRi0kt3kkb7JsrVNE7dpcbwqkp8FjL9DuqtlhW0PpzBHJYqXgL138xBUMv/efMeqXHlK+2KsmhNA
EqeS2UO6qNJsV9XMK6vNsT0KjJfDnbaSjs/fif7UFgUrPJ22lPHs+r0wNGDdnCvl3hEbvvmx5mQk
dxAEAdERKMPnbJfSRRZkQ7aEnQEwQNFGdDWYP/ak4sXuzQGcn5UbYhyWWiSfnIH1/xp0TzEqWa0z
+tMdx63XY+zKNGnPioCHN0VhQ7m6igM55/NDvkhxfdVeS0SN1jaHflJp9lXViYB+FdEvHoysgxrt
Ii+ZGhxxc5cBXkupe3mV5e4X8fPHjkyKA8v90w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4208)
`protect data_block
uLkgvFlhr3142315Ki7dD1iBKaQMl27DPqjt2S1iIXLKlbU0TdNHdBx3C36kB6Lhvz41cnD7yuLe
nu4U27rkaHsVNDPsTVJ2wsNYxpUCCOgMCtbfiXS8K7hEKm6CSHalP5/9P1CNciiOYr3IKz0GG99y
0Fm6n+0c8y2g3OHgznqrxFaqC8jTK0uXRm18cBlwPgp83axtM5hQmO/AeQnBNA1C97VaSHBbGZKx
j4pQxozvUBummxnHJXx973FZ1krNfngAKYMcurW6KTVNq6TcqPImOKxBjdlYBLl+IALpZHbc0IEY
BbHmi7SIiNgLFfen51zpLfPws7ZZKo3KRKuvPy8ubhS/0cjasK5ji+eZxYaNQLf9fwtBf2W4/FaD
FCowbFJz87xNlLT+/NKtGl07wjlSw/311vY91/jU6nTRPB3wqwz0AdOhiNYpkCq9FOJclbS+7+/P
N4nit8djjYvHjMndGkfXVXfrI072V96SM5DzOX+1FRGlIcVl1S2IbIdzjvx9XCMM/8SHIBWnDT6b
o0mKlV3dOLfhAJTDZCE2rfIjfRPCQyIxY8+T+j1hhkhjenaN8zRWHykh4W/p7cBLy8gKFYKqvDr0
AEHeq4ZXmHcV/OIqRzL0TDK6ZK1D0qySkJ5ZeK5hyVKdYjo+/nYsCAULeHZbf2Zrg9rOIbH69/Gu
Y7esL1wkWCihmOCqfwN4MlYAstpJ6Mx0w/Np/pEaR6LWNnW3zdQ3AWGYeHEN7uC/zyf1D/o0ShbN
rzSDejtOGqDxTgxKKhvqBAi6rOKQEgbqGizCVT6axPZztwZQcrCZcpABngf9EygZ9OB8w+IMxM0t
tBkhO7R6ojLgK6TECu4L4P0HXSr+PCwPuYA5MTlbZqmM05EWLWmsFdGqAt/U9woGyfESCPnDc16L
a5XmPpJoawfOcpHRg1+DSwUdX9UFmD9rTHkG6LLQBIUK0sZZib5/VfGi5A87naQoqvflbNLdWDjI
InbE8YpXQ1ACJpEMUT34b9f3DRIlPIdhYsBXCJhbc27iwtErclLEZlcduFTcH+M7GkSVmakWlzIF
euZCo8ooQjsB94BobkmJtXG3ecIo2h5ycjTj0Ef5PJGVWA7KH4g17FxwkL/CJ+Poq4aFOFZtwvlk
FTqxee9wU68TTQPVUVer0zccNJlhN+VB6USU4x/BiOBRcUD9P7HjvP9UFq795x6CYHT4NcJ4joUx
mJJ30wGAScqirQmOnhdvBf6nnvDSXwNYWLu6Hnt/Q484b8LpgZJQTOrWIljen38IVbg90QhUYRyV
6CJZxonQzDiZ3wkShRq1CdI8NLqqEiUqSHKs/EpRMJYSPy1bb5/O27X/XRNTYiQjutXGr6904a3f
yf0GiWo4+1xSwHvMNj0ECDgpLja/HRRr9yy0Shs1EnF64UFQOKgDgXWPI8Srr539qCLWmN2P4QJR
Bn231wnoWEL+wzuBJ69DJ75iOetv+2MYW1muOffKwA1E5hxYVi2rTVppVKDPmAAWIXvAXck/oIOg
IsgIqNY6Z5hvFr9ZZA/Y/C8u1V+xHbGJ/9+zarOquoonJaAsZN+Lmh+muvVx8dY+ZCvsrje4D97N
6sjNm84MbDAgsfn8MvLuIU02hdH6cCy89bfonCaQs4r8oKHIZoII37uCW3E9Zmdca2v5CeBrl25q
wXhXmJ/vC38ngd20LvjHLxojl+xRsbcT4WpWGP1fS3NhTggTSnKUvybkJ9lMA+uSv1J88cdyuKK2
i3VnF6PjwsPZra3vusngrcavk1UnMQPCz8NBTy3AQ42/uIvZli+fmlEr3QCSWrWdpHFEVC9bUjvm
Ozp6briLC2w7qe9VEpUA4EfvadpAK2OtSYfFNUIDtUwvpqgVrQ1SAln4nhGQtbWgdaJqdc3PzlCR
Bkb3ZPoA+09Us10hIV/Z68y81eJMvegdOFPSel5GvwOQADSKbsUGYTn5yKP7ZByrGIK7teoTZMT7
i/5+jCMW65c153hD2J55w8ZyePSHu0ni3rIl7qVGy3wfLEjxZDEAeQC2j7TZHXyVb6I4teDPgrc0
UX1i1PHAexViI9kWkprJntA/+SU1kXmfMbSzW6EmQzyzQ/TejASVf1+OcpFYrlzC02Bp3gmR2UZf
fhU4YtGkq/69c3T4OshBfkWRHWqm7Ko2In4+OVjyEMkq6zqTXa6NxH1aELeZvb95fEeL3sBBerl5
arS6TRZl1l1sNh3Aclvu7wAGOzWcyJbAXGRoBRqgVOpRYmUVrpCpg6BGJ3jrZewnO7+BoIOw4MKK
A6U3CnXfgahTaZyCUYWpRFRPd+nYmuDKwGn55DYsOFen5NKSDF5dhFIUb813lgrMGIIo99Z6FAEB
bvz+v+3g5CPOjj07alnIphdsPQFwjsl2BLpJs9XhRBfPS90IVmOPmaXp26Rg++l0yM8XHenA/ZUb
PKsrUAv+8C3B1w7hGT30dgLQ5taxTrQ+6lZ4yOzda6J3K6LhC372+Imvss+HGb8SAJKTPS9Vi+jZ
y555d9lgUGh4EqruLQtanN1pFR8UOsbXr1MBQuPt0wijOWEGyfyfc/IsgbZ/QJLWXEkLo5C1X+vv
4xxY3nBYu6uXJ4WKtkHXeRn1Q7jRQNU85kvjmpxuovg68tFXry/uGJmR9Bs16+WNgbQ4jLrw6frF
DlMqYnbxkr9rN2A4SQbfaIU5+wNOGcXcwJ15fIHTC5+32VuP3SJL8+NCAOu/vrWVLuYDsVrl4mEP
3hj+iDfdJ2p2ekcLHESbc4ETCJiJJyue5v+cWpcqU5Lx140dL9c30GJ4EFfeL6qoAeSyCSG+Z3o+
0p5v0yNJoSMkalXoGlfpjP1eCnV6Ww+352km9OinVk0En3nkHaC1bj7rYtJAlomeJPoIbBHWlmjn
iz/UUXdZ3Oy0ggqNlZ4+GQvhVKoB2tCNVDMB1wwxdKu9eslzJrP85KMsamppVi0ratGmcWKiluz8
WOp1Q70NdQlCGit3b/v4Z1xK6k1v0lnjviyCWhd1pevYysRKTM7h4Ei2GeEcXtA0k57aouVaZxpR
5W5mObf2StW9kAbVzdjA22xHFbBD9Y7tVpH6cQdzrX3X3e0woVOtyoqO8CEnVQNxVkPBg3kYu+2a
xroYnvoWxu8uNCKBBpV3nD0xtjnDrQiC6kfjhUJZ3bzA6OCZjWqH4KvD5Xc9HZ8rbNKR5elbXiDC
4Fx0IbZTPnlwDHpQ4Dsq7kL5enp6ATGcNeJTqtI5VmzylB67IEAKN3SNBcRDYky7ul5XP4pzpmtJ
1QZEjd4vnqqYdJ7bsGDqWueNCgaPGwcMKi074z0zPp2mzcxFlJovzea7lJQtX0V0ILlH928cEuN6
RMPR63SMEOtBTc8Ry57gALKnETfmjvv5WLpw0H8DRdkQ2Z8na/Ol9X8hg+8QbEexlnkW41iGh3aX
NKR3NZZXd3YZf0ZIZdalMf+c0vEXAb914w0SAzXkZlnRE+piZVHf614LsLv23CF43NYYCWmmauu9
hWMGyd1smVBix7L5wXZVPOj6K5TipqpXA8HVRE3Yjgi8LzsZFysp0g67pYt+BBtY28h63tOfS0DL
1jqpwLdouaa3xgmIu09zC2N6aG3iB2C5J1MEl7e6RK1oIFLYlvgFqvvR0Q8GaQ2NSGG+qNTHIWpP
5n1MhoFE/EKL1EyJSy1iJyY8TGhw2VUBoolU9DvJXZUTFUcmot0Inf6Yk6PD1dV3k5zoW+6fdhs1
gGCsy4pcD1epiSHRGBLiGfNHJYd5ZkuzVrts5v7e5C68njoz3lD7b2msXRW2I8Gz8/gm+/3ISHIj
7xmCeY1lMue6g78lFCP4fX+5dyGMy7qt79uJnIMQnBzFDOh2eCMWdiYp36LdNYAQZksPb+pVfhtH
+IOPTIvP0JeOJ7GMKpZc4DzWYdUtd8wuHpqPFgYqLoOVPyGN87ugXapvfC2Xzbp6oOgSI631nmem
tFIYk+o+Q0jo9UeWbxelzlPut2LsWYWRz8b5PozWputxzoyuUO/p3+XZY5KwaY4uad/P9EKmYbXr
qxAE3JAMt8P4N6TEzYinCORgJHR4MKK8v96d4d4fXk79VY1N40NOEbWYh8BL0zaA6QsUsDu9SoGB
Rh24NEuS0Im04BTqaV7bMb8i5gRfErDDazTPZcPl7XybHKc4coQYerH6I6Egn8HlPx36bZkg64fd
AwJfFcxDPDzy+INr23JUclZGdfRXhe7o4tauF0Ss6sy9s06ZlubO3I/PfaVNFA3cp/Q3HDVeASFG
zhSQ9gR9mCpm+A1TzX9roZYbq6jlFy4FmxZ3kKlC4jdJOo+Kb9nXvRMpinNNwGzmKSwXwASNMsLc
/ghk3KyMIknTWBiRO3vcQd8AhPZmUrhBTYiYDnYELrfq03clClIhzLz4B+VhRIgqsoYd/xW/vGxh
oBDzG9tgyBYAcO7FreaQR+KAPUZRt4z5FH+wpObPG+c/M7B33JamxeCWaV5hW7w5hKUj3pRlkEqi
DxzgURWUoWAHxMuZ4Mf2TjI4ogvnZffJ2HfQjh/VqpYj0lXcwhesmxxIfS3E1JW1YSJjxVl8WlaU
we2IF1KvVxl+hGIfhrY6EItIfm5xx3hwEkHXD3z2jynjeeUEzg4dI5VfBAkRfesKk4ZE4+YpEj8w
sdVV4PVF6GhokQiogazc01sm27lYK21O0cJql5mThwe65DyAq8GS2oY7MlCKQz6imXTTPVWL4ZOH
4xAOlCCF+Ig5WieJwSfjgUsFE4ZdomsasNhOhcqVW8LUXgkNgjDhzifUB6mUF84HTbXsjvVHERq1
Sm2gFDKEXZIH6PUFw39hEKTVXPwXVVjnodiESxSfNN2hNzIk05iIbvf0aGw+E+Hroo0l3F10/rvJ
eKljFYU2vz3n76+Da796QO7Q997JANUIZsS8n+Ar+yMzj2j8yZBatRDEAIgIXZjD8R+sOc1otWfI
NmoOrPRvE1v9eeGDDloKBWBodsserztyBj8AXFc9ZfBylz3sGDwfHkqcTtm0g1oxBxxVkdBQplsz
2D8CnNbdonQCUg/YeySk2RjzMu7+QNkIYt7sZlK+GsE3jFSxu5plNRdhMDjtXWD1MEEkiHKcABmF
ooLju2d5ZUYCkj3WH5ir44sadBpqN9D6D0s7uLLWL9YYrHgvJu1prC0FYpV4HdgoT+CFKmV6Kbwp
PgyCXkeOIbXZ2Vb+eT6gyB7AXFUJrbp06jt3XQ3LFJpyuYL+uZQmQGpYOrESMIVkhjPI3ofH0/2b
ZJi6oJSsujCfU2LnuhGwg72BVwW/pHmf+yuvn7EaogS0wmwoVB+3fSs1fjKljcmTvA/An94tPoMK
c3yAcfdRYHx47xrTAHHC0SzmJNuxyhD6RWdEWxb+MJjhs127rX8kxjP23+HEEWMAzU6rOnhakaz3
LekVSqfJ+I5J6LMu0QgzxohPaJPGYXIb8iE6d1yohmlcndDa50MhonU3dYz13seNBq1IRmjOSCgG
Ww6OCWZRbx2doYeFVBJ6a7c/EQQzCLc873upYZEIfAzQEv55ukqZEEzdev+W55uqC+m/SDW5rbJu
+ounmJj/mVnD2Z+/S6fFaZN4rGW8hlmzKtMHOtAtBNehdtey2hDkKZ+YMJNZlJY=
`protect end_protected
