-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
NRBOt6jgKpk5iGHiZHdABLlyvLLlwhZUGRllNSci8FafplKpe5+odoBefVtwLo8cbIcfiPOAzFa+
HiAgqjpMkyoSCfbsNA9Az5Xs4uVSaUZbBTlRsPLjOUie0Mvudqp/tmxkoB6/Ryz4qiL7sZa9cIYe
1jFzokleIeDw4BiQq72GcQDgm8jeuPOiGKiKwazBq0hegCC/2Qesae2nqKtNisd0SFmbRa0Mn3Xl
kCiNqkdEkRD0lJw910C6SFCvGINRsIjv1NFqhkMyLKkHxZ1EXlT91dUy8Z9F6LF6G2N1HffJy7O2
6w7UpITpGrkU4N7XAmDtRHrmKSmpntwzKEjbjA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 21232)
`protect data_block
NwFtmm0jLhMfh8M0sFMmY7IQfvjpa+lrqFqNhXcxjFu39H470TIkmciEXc6VR3a1FW+jaHys5iHv
XBm0JAP/6nVrfOEaH8bXOhUHuLvEkunFdN9T8F6BIRy+59IDapH3R/GtETLIdh4QjkgpJGNA58P1
/PFw3zxgPF9j0D34uI0i45uz5ePXudvuZBOP0yNUSjJuZ65zJV5roihfpG0SrIGEfYZLkdsa+txZ
g3Uf9Bmg/NDSL7fCxfJIo54i3MEa2HeC4oCzJg+eUgxxjJGk5vwJHehZ4qtAVKYl56H8S5N2BH/Y
1LmQeh0OagDDrg/fwVrFCK13GFmcednO87CepoowxfOP0ebHFsSEx4xjaiYdqT+48CzLZZvkNgWi
prnOAUk0qynYYmiQrfo5cJYeu5PTT9BskE/3+9TWodIeTyY6t0Ue89Ixs2EgDt+61m4XsXCEz5fk
98TurCN+9lz3onfeAKw9o5iuDJvwbRNOIxCAZUCTbBfcqf4c+HBi24wpjZdHpeitXJkQ79E2lvFD
5y8LxNazPqwtCm7GgFNZtpH+OAIiEtTe0r2q4uyd21HZGAz7cw62wgCANAuju9aJp00S74Agru5V
0+QPZ27TbCZQIJ3TCb1dNZj7LA4jLmJgqQ6WgrgJJ0XyxnCUwOytxlilBxlmQ6Yu5zt6gMMDm8xk
hfI0r7CO4sUF3qBNydnguCbCC0CK9QHO0CqZn5RHRDL7R4EL3B3jzzfUykApzVaPqvhgNBaxHiU3
z90dgdXA7CFJ0UnJBYjz5GimPLDuoSLxJFbyzxRFd9nQHObhkC4Dzu6EKF8jA3hPL/3SULaZXnek
Ga7/g7BTGMkz5p6VaPR+QW+ORgDH2jaGaWSS4+P39ET7Oan3QqSSLw2ODq25ED7HVNTSU9hpbyZZ
ljmyQefdfUmS9ThlKBtQrUZplX7s15HZzDN26O1NKnUiiEVFmdyJuQiFkQ/hZYJtG9c1th7pxQeN
qx8hmed7Kr2PQcPamkyEhDi5tq1ajUrd871Davct54lCSNMeyneceM7YlmuhWO1Yir1YQkSndska
4CQ72Elrn9TSDSv7gfEwOTTI2HTFGGURyDcuoD/3faCsAfUMMBNb2EZnUjcYu5IqJaen3dNjbToq
aK2tTcxOOMz16C8OFt0/ISlDROdkMdoFg7tN89Xjt8LoqWnFhOqIQLhiarzYa1e4JdjOnJskLhxT
o3oHsd0sejU9wqu89HXHE9bEu3at4nflol6UXtv64Fkt/SwEd7qW/x33XRvYMQP79Ks9tsp75oF6
bYAEYlCAViwyomo9VhLDGBznnhHX7K6IpJAGB6coEYij1iQn60XB215gGtjO/U28DXqRulXkrrJ2
T4noRRJwmipzEcc1eB/PEji6/oZTh5rwhskshWutwBSsUGQ4olh+8mIrvzvAFmD6RH8MhGwxzbVf
ryO/RaTaQY5b3nCFbvfR0Y1YpMyubg8hQBPm/go24f3wWEPd1f7IZZohkjhdnD22roNF2EcSmorp
Rctfa5j08RR1g7y3GI7xrODvxT0tr5HpdJ/rNOjKb3WfjkcVCCsJmkDufpmoO/5zcn5xh4WluTGe
vt/d2AXxhgpctjH2JRmhCBpsi1nm68gCkD4Z3OxYcktFNn0iPnKuVgjATsh+wpu4urRITeQQTFvW
il2TD2Ouga0bjMeVAPzu6POXl+2erYOp+NvGU+czVqj6zJtNfjJW9tvlO+5GFPgd68LaxaqlcJr9
4vXfPbnUm+J9d5E14E3bRajdHnktiqloSRSsWG5CPh7KF+nbF96Lg/T5mvMVCRMzN1ry5QErEjaJ
wJQFtl5x1mbyvBmWB0NOZuY+6EkwUP+qr5ce2f5xezTohKXZnW9u4fbUvLqEml++wdNknPeI7R4q
miG88l3tl9UWjqUFYD8V+NtvUo0C4lM4STrKeKrWgyFTIz3rsiXA6T9phbf6zUXTLjBNfKorrZbg
N5Gt3SVqU4G+0P7mEao4AAyMHUNr2bfqpk8hkHkUOTpLBtZr+MED5zgUeGV+iqIgXpMhfwcxnvtp
fRCkuQ0bYUQCuPtcoZGooueM8HHzGMvMDv7RVh7mSnijt2fZl5860P0m0cqCthVq4Oq+3VqfuibT
MK2VlnmQJ7IiNK4Cdz+//cyHn+nwz8ijEjTkbGpjIrtPGJryW1k374S82ioqLFVOld3N4kLbq6Jb
kVGDRGGXMkK7nxFZJEI4m9hEDawWYxFaR69DTAOaeGwrfojGwWEbeSUKsQ6CVOztgls7gZ1B5LUd
HAynxORgd10ncZwngsTySwsnzbt6fSjyMMKDDqlvILAHmUnNARS6Ut8pAvgmJMr7EIa7QSElVJ4S
ZKkFTV3DkbVzgzPszXHAqTp3v4nfWLrVnH+Gy490Fa/Cz6FZDg7wl5b+CXQzCp+qlaH5OeZpOcX+
O3D/fVyXZOLm66Fg3xonfkwUKpSziaAzf10F1tKGuOM6BgpDLgPrNqQgc2I4k9MuCCxONSHs64LR
P5xU7PUW3my8MsHWtsOewEFT82bDm8nIod8pJb9lLP48MAUgvKiZyKN33p9ksG7KZLU3pLxVqZeq
SsknEqARNVnpfk8UXXF0kBa5XZOjt5mkj0/KTQQneuW8KEVhIvcKqW6DkeV3RY57voXlhwUSp12G
qN4aqtXkH3HDg249e4AoLBpPvFOp/NoX9FrUBgPcavn8DY9dOEx8v5ZNDF/gwz2jFeXhOwSr81fe
A7ZaGgBsZr+ZoRFCWiHTkwsFgfraSwdCnuaZlkHMXPCMSBjfkzJ7EaP6Ey11TVsFB3Q+o8uXIWjr
BQesz08OtRadfeGdfD2EbVUx7liR8u3ziqjQDRf+07jzCXpOxPizuqH/sOZv/9F5r2n/rQhGf22L
dapvbTCNCwHR5IdwdMZU/p9j8+eXiwfaee1BBL/PzPNv0EdDjtf7WILrtL1rmuDLIqwKWigNath1
pVoz4v8xUr1VLwLKSoFj1q/fcKB8+xh7TJCpDkit4NOcw4wvlzEK8UZdFXl9ZNK2gEDpGHg29l6I
b9+ibDIhIlN76Xu7ubkbGKrbEUhji8kJ7LLpTOEE1RXFF7xPDg2oQnPsspcJqVv45DYtDekm5Bk4
K5qbHuJ2gZF13CixbMIMZo06dUtauthAU5MSM8M/XQyjLWDXqrHYm6dgM+uBxT9Vq7MiphOHhsRZ
PGAgGzbeY8Zx++zEfHSIUTcIX07YFhyjfgQ/9UPC/iKm6AWca9qE4hGuKJha0RYeoUQ+WGAMt5Oy
20I/HF+vovYXaDx39Z+RKiebhvNhSy3Cx2UP2PuuUj/witxl9+eF60SfijH0PJsksZzCK2uMQlo5
kvBQYVFoy8P2T13g447H7uAhv5tQjSYHWZlhjDMzu3HjQNvUAjHTmTfszxn1syeXib/nHMsxQnKW
9Gycn7dMVVf2AX+x2NFZuOKhKSekkV0v0tTb0xudQaa+187w+/bWQS8MK4GjWlJYQRDuS7OH2K+8
aY7JGXWa/rwMkmKaJwn/Jz5u2gUnDLDzFQpy16ECTM9JlmNTwVtI3g2K/9x/M/TkYT74DOrd20Fn
mdscua2kYmBU+JikQwCE483MJRIFRzSp6rAiyzKcS9a/F4wcSw9/vQqD1e1qkKRaM8QHZ8bwFqQn
j5WjpzdJQOqjITkC64jMiwrTKgx9BKJD2ZaFzQbIhtu0J15egSxVLCRVr+s2MwuRorKJr61SHKy5
MEI+3yuZYNC3bjQirytVRtEBDasYwdkB3tcd32hETiLsa412wh8MTQ/THdZ/lC1GIDRrYivavM6i
Il86apMrXG1yPVVRHTzuISZbCd7VVerjGnqP7BglIy8GiSg8QJXhc2xDIViORhYsQMrGindVpyA+
iEq7bF4QPvTvZFFl18LnJmYJCw4Fh/WMMkn2luR+6V9OJlGAHWRltciLYfTg8LZcS3wSedSZHqtL
fU0lIPpznSxiGjmkPb9s6uWs8T/4cYzloKZtIDSLv7CIa5AQNVJOQ1AwUK8sUTHP5N8IlhPRKkcB
Gl0lO+gpvO4pWW1OIHCLFUG2opW/yJoiov7yYJ4nPifV9xTPNwy9J945TTnHrjFtJuV+jSfhtRVw
BJQkRvGbDfUkDw4K5ZUGmO0sCB8sVXGwasBMym/i/C6Xi89wjOUcc+A1oB49pQ9tfRigCr9bWXpN
DqXfgh6+FQE0XsOpV/t3bj9SB55ejyorAAI+4jjXt2+qqdvTrcrK0R0dzLUmEI9fSmorEXpoRlNe
nqpXAK2aB2ODQ2M39YcYe8ouZJOBkw+XnfdVb8hrxygiIcRVoiioMyXBT6KPx4+PZeERGEsp1MpQ
L9hPIZYRIQ9AZI3sHEO3IRUTfNHRK73PYyfQQ0Qk88fJHWkqHrr9j2zpeo0/g+L7EuXgmX8qJjub
gwmOfEFal0Gj4AbS7EC8fLiyPeuEftfHgxpSk7gu7J/FshVP73lT8rIlDxyiYBF6BOZgzJ0PC43K
TqMkYKt9DAP3+Vu9hADl9d0ulZKJSw81Oo8O4o6O+RoJTwGQFeFnmBVAWo7jEDMYeys/WL7+KMse
HSKv8lJ7is5t69Nf3vrAyifZHGdafRo4ZY8yRR7OU9zDFat+wqDc7OEu6zQk5Kw42baq6E8ZhtuW
z0bEJz7SQuzx7WjmywdGwZ3uxPtEITQY5BDrW5uDA4G8Mvip6+Um0cWpXiggfBGmCDyWmRO9RjF1
Nu2igHQW3RfG/5CuTqSxWL1p5xwD51rb1d6jGxS+TdSq/X2r+FDZmf2SzdPj4yLSvSPaRSHDsDf9
4/0OjCA+D401n+Lj1TX1liY2ZU9iSbCjip++PpYOgJi6hbsoTGO1XCu+LRgIM0gWkzzbTbpE7GEd
4gnf+CtHQJbBPGaphkS1YaoMVDOb7HRmIPqUtQf9GmMSnOZDyJ+Lynp0hidghFK65+qXgR+dKrkv
IH0QnqEDT59DF8MSlBMW9+qlHL2r4V1u+kYK13iGcsNSIbOMNtqORWVcq867sr0I67nFaEPwdZBu
WoNX2CmhOXgMDdiwepTUj7KNI67ECcG8Tyh8WfdgKBMhTMwKgZLod0rpOcha+yTtxAoYFlL/vnbT
txiG75QG0UmdWNHd9307iwczVOEw7/szxMuVnonfTLZj1M9mA32f4q1j+X2M+JrAzWyBCGDpIZmt
8QHrdqZZySs4ZcdMOvF33uW3NDsrI4VpgGiUljvauvIaYhTlQuicFAPXRIxBGKLBalfpGWwbGm9g
oYRo9L3UYaTTSEagebLQ+i8cNOvAM49Q78qtpHOk1/INM77EYf4tKP1REwpp/B27B3cET/rUoEoK
KbHTOWdJ/A3Efs3i583gti5UISBnb/XVweSTrLaxrwopow4Dte0Le6z4o4U/1YD1s2YbCFU8SD1S
tEVOygxcCM9b8ETjznQewbJEW9Amkw47qTf+9WLIBFODZ5F4+F9TqT/tKobwJomoVy19+jyissn1
SNkwnxb2OXCjQB2MEubBA+GEifUciy7LEimPK6a3vWVJaQP56T7fFJOUqAiuD628DBPsnFiuVl0R
YiaSogqGxhC6rwlQBY5ARi1iRGs8JwhDjvnDqYbKx8EavWTiyvGjbGvlUHElfZyjzVINvtcOf+o1
1TOXb5bNzbTecJpwxWL+p6qJTPQFHyaWdZuX7DJQ+0nCkvct8aC7fck9X9dXEK18Mf6ojlpMAIYV
zdg6P8c66PBzRyiV+Qlxa4X9aDgLS60Pho3oc4Jr4PSgTRWZaFp5dNpH2gQzYKRJ9C2LizGiewPC
Nsune4F+q+PgP6btbtZDjtmE94N/stoGIXJ5ptL4iBXjDN92PCibgFksgt5DJfccHRjwsE/gYsY7
BDRS+xZxblkrngC05K3Pt3yVEshCS8qtBmk3fq0yT+dN07G3JyxazzJbR02yCKuVn1F02CMrRWTF
XcacI8hl46xblM8xMxvYe2XavQ1Tk5lTPzt2vu1S7uwLAt7SlUJpYpXtmx10v8XWW0XMG/2I0mNn
vkEfZ+maC9sWyN8aQ8f4t9F6O9XxXG8tvjJ4ZuuYbcUQhT9JO3wJXdyogYeAzMB6cr3Bn8ay+8LH
OCKB9EZ1wm7hgoF/23vWTKS6lGWE/CoWi04WK1J6/mclEEFQshDyYoW4anBCR2NHjTBOurswuCPH
SSMhRMAG0iNChbwIW9zVMfHmhcZj5vq3s+nBVkhWMNwdvmse7669mHqU9u1KmUy5nDOKyhfZ5we9
WsrPefyFuzg0S6zp5/86AR14CIwrAEC1WMVSaXAkE3wKGS0OiluF+TyE46sGQKsvTgsRmOWHHunp
nsHm1g/lmzhkSi9BHf6m8g+YB+fIUQjLSVERHJ33TW0GcaMZPz0FdGrDEsEyOqy2uYwJIwA1b3n6
SjH1BxmVQLIYHkStGCAhxZK7vlr1eBWP2nMXL2cCPcHwArHvatJ+3erL4nGPfC8I5243SPP3mYGA
0VRb209/1XmFsViGHUYeBsb7TTuW+Uf++ZxusEdeFQR5PSIKGA4DtXTnm/BMV4C7aCWennMCDykA
D7S82gBzy2bq4rtCqKHdSwgYk/IbzHGu3dfmu7svC3aDmRLehVBzMqpPp4bwsplCUnzdGrpRVGJl
etYsfYnbMFOqcTYcfdXpj7lV/l0IlA9ImNF9dFijO1PiYbehCCocYjrmwHwCxD2Upo8g5KvsPFUO
TpZo8qFgzcvjIqRUAy64ZDBN6IFmia1KZ+s1gCzRInznkuTclJ2+YLLAqxMn04MtiLFQPCFw4eF5
4M8AT2+SRyURoB86G6l5tbMkW3Whpn/812+e8+G1+HC8D3BGS4RhJS/PKHtSLj4nYlvVGeKibi26
jivRE827ok2b3C57mXVD5IKWzAvFyWoPboJP9nDGT0g9bv8skePOXqkG7znRcWrzQullJJsRh1vp
5/1TRBH6Ls/lP8Tv8quSYD/8AqZf76a56wWheKxkCZ9vV915BOPor2/2MvrYJKCjygoml4huWZX/
zno6kwAK8aLjKBNCMuBezV5m5Kq2wBIjXMScsOK+fdyaLSxpXwLjoEIHWRnHn8RHiZ3MZ0wnswkL
9EOU2t0qp0kVxJ/lmeMKF62uWmbzelN9ure4qnW7NxXzlEmxFJcSZmppdsYyM8RbPIvsO1Fs/qn1
VfjqF9y20M2Czia5/DTcBMhw0axLPWq9IqSS4fcT32uNGdRKnb41aVpf94wISuZVF+jwpzCyNIJY
nD2jY92L5qWk4Lo8Q//9eypBOgkcJb/Vlng+Q+och25zxqowFLjPFXUzkzh16RJYZXphXSPA5Ut2
FEUn9X3l9m4WTlFt4OPDKvJQ8HLNMAxWdeZOrHke15FaZKltO1h6gg4Uegb8MxaDBJeOzd0ICdcw
Luk0kRfMJbr0/pq0QCxvNUwAzkUCjcTimUxu09HvLj7HqOW5Wzn253Xg8MEPWT7FD9y9x5pY3nzF
RKH9wm6EI9XbgIRgG3Fv2C6MELySVlL8kJwoBcj+qL5fONCiua3p7uu0XiRs61pODRxuMHxfM9AG
V5xrPCJQT15aF/WJmDWj7zWA6OH/HjnXR0B7FxlCl/ekNc0YtlY8rdoNPfwOglxhchOjnGrX84bZ
Z3DaDaNXtucswAr3WcyxT5xbFFqcx2CcyIxx3zRJ/mOIfahU9NagdsQDrV+rFRCrt+aMlm+o/G7H
sP67cOMDn8W45rJzsavx7FM+xtpIGc0e/UhhyKVOZUZ7rwH+NHiTtCMG7gVYh4Ihv5vf2143ZFBG
KcOFFHp7ql4jOGz99Cedf2NxijETUWNpBBu5qSirXkwiBk2Pow0HEZQRdyNCAe/Zm7KWnZADyp5u
pCTBoBfeg8OlRIFmMDZzEKyh89yn48yW4YcmEIoN/8kwCSREmt/FZTC1sV8dJvKY8nnJ2PX1uvLl
Lj4oEFdGUpKqVee4ff2EP5nwFZBzin3K1Adt+8ysLovsz5Rk5xZ9pYJTDDELVCq9Cv0F+uFs9WQf
aAWrtAuyv+lGCkVCJ461P4FDgon/MP665rffR9mZttBOgU4J0ZBsErMB/BgUFDNKrc3VRRJcTXGb
MotpSmOfNch0iLeP+PE1ye1Ryra1nVANeqF4+kY5ciRuUC+jRWaEDsTMifwzv8JDmx9yF4kNb13S
FxmjEFf3HeaEzBffBDqhRZyFnWKfZmrO4xXM8ZAwiAni58TI9QDRf6W9XMOZTi1dmHyvhmcjeyiR
I55QQo84lR52qJNwTJ5DHq4uiodTv9OnYXF/ygQGKgOZw8wwwEd3WULYjgNRI5JcLJiA7bwsKHR7
FO3fvk12Ve4WoIfS9c1YLXe2gBFxos5CjCshx4wgyi6l+hsqJTM3zvI2hktkpd6xVDxoIDTOB/YR
cuVi1n5KWjnghWPxflJDQdpd8SiowJsg36zhKpDXVuXioxjZzEvjQuzNvED+FZ6iOTs9YFIwcuMY
X8PwmB61EQXgUlDLTB5kJctMII4aPqx3rVQ0N8XTWt7i/B7w4XSgNSMqu7tCPMrxo6PKWEhQl+BX
oM/DMQ4adKRMKj+76dseewPmb6XWjq3frcKQiRJBrP224GTUXNDf227uw7CfgK5gije6B0hIXK7B
Ei35OYW8h1KKjNdL9pYinSEia5xp/wgqmt5/7gK2aMXdgJFTGklgcukdHyoZvwfj23v9ZTJbmhDs
sgNKJdfHQs5uQxI94tN7gADmwEJy8F/gn4hd+0pT0U4Sq3ewHhM8P8dAY2XhbWlNevUjorzr9qQS
dYGbgoIpX4ODe3bcChla08ENx9nrSc8obFKEcA181O6ZOL3F5M5tSapwYPPJMBB6JC/pXQyxVdmQ
H1p7SFNOH1c4eZKNO6CEVBvdXIGKV9bBYrgCK8q4rwp1MIdEOvFwiDGrdE+RIq5TsbQY8FpIuP0Z
SCYecsPsB/9l8HDZrUm+3Rj2Dgzwwx9pkO3eafGSmY95TYB23UrzRpacedBABRvtlzPeS7JyDK25
w2H9Zj9/MCXrtRNxHCNasc4FIsbQOcP5JdaSDJdYR7ewU4gZcqenkEtWeALq+7SvgQ5bWnXZxT8j
dUMnZtXBCgTmFMZkiVH0Fvqk6ZnQ6gXqCUw3r6Flt/JHyYrw6UiuD8307vphxPZzM5ZkB+unblBD
QO1IhkfQCZ10WwrL6bPoaCSbuswX1KSIZ8trqjNQAAGHbjP+q1WSRsA8TYdUoET3DHGbVVa5lbqA
kKIA5M+PWRUkpzODN37qLUh0umGrFf81/k20jFyjOgWNBa1/IZqqeI/JYwXaN2Zf3WvY+o88waTe
/3PStAC/BhAO1g+MFfI0m1+tMi+sfInz6qx7AkG7DMToLPiZx1bD5n/GDjr5jRwmhnYGlgIasaQM
MZtG5+m1GqGhw9+Mx91nLslfxLHkooaiKwBPP3j/NnnswqwHxMDisVyG5fs6NUxs7aN0xZ8+/nfe
a9CdTwTO0E8VKTexgULRonp8cfOaAjpdurQnmQmmioj0WZ2fC84BWfTNfQ1PGoeDOcu4+QzRXPQa
sTrSXwtxI9gWzhUFIGiI1FHOvyKxxuU9QMrDT//mC/OisZLIag4liWyKbkgzkVpAMwX8JVd9atM7
kIVS8nNDOPOzTJ//rYSR9RGMZjaAD3Y4MctklE5CSAi0lnuDX3KoixCSwXjcw40unpptoOvgpJha
WPrK9CesKLUhIjVajlpJ0fHAppVs9yscF1GzPahXPPK4tflda1i99VXp+gftZC9MSoVWyCpjabY+
KWwlM34q1sIAg7biekftTUz70ZEHHOjlGLPy3ptfR6OnXvKeIad0PN3eUToOwxU3RomY4a4kZtlo
2Cc4lx2g5I6gqHEkS4qUPj5/nyjm2btUnQWMfC2AazRHSNEE2h2pAGqCukjHtBhZwou9u7joGNVx
aPIZG9YhgXnX9B9HqzvB32SS0dPN1c0hqSWo1bya8Pl1EBWk2ku23mF9ud5JghGuIgDZCm56b0Nd
CoK65GgysVWoNybhp9/D52IqPRf1wBW2PCf/VtvS8N835k0RX0hhMCwH+5lqWhtFof4GSTgt7W/g
yjJTNw2rUK+PFHcQZH1hlZ2M1Wb7It5gGyECzmCqWB4DgMH6chbSCKZc2WeNxSp6J16Oyz6HDGeq
JfBqA++1AsU/nrhTpaySsLe2zc2zfvi0yPKAuRM8o5LDk60hgy5HcN0+PfaH5ILxd1SzELusRACV
11Ou3m9xgqRey2GpG/JKnRB71VNUyyuy9HEJLfq4pnrmG8XPTkPoTRC2ezjc4JYaoHO+4iA3Q35H
k8empCjuzOIsi8xeF/vOYJ7pukDCan4OQ4uzO/98/OD6qk3MnmwVGOOqBvsClBEAfxh0P+vCnCtz
GxZ6B/vcOJo93Z2/P8GHVIIkKYHP9hSwTBIqWTn0zAam9ib7nfb9h9AkaUjOjdmO0XCVZxiklY75
VHEkh7Kv5CgwvQWGXF0YMmJDTrLbNHc3bnf96LmzdTwuee962rOfGjTmdR6E0VH1qwK02d9I4acN
sfGhwstjDLv0jq7H22X0SASYsbOPr5lyyGyHiGJJYHeKyk72O3VweJ15BbOlZUDbkZ3ZLdjGYxlA
n8tNiq32HDnvjhhKzcLEN3Vm/RonzbJLUHamRWuj8EBk8csyri3iuO3gE93PJGaZBX1zWWwpIwfK
8JJr25tOnpbFQx3vOWDM6Ati1TXvt/yN3IhsA0x3autw5112IuNtGJ4756lYOsq1aCQKkzrybKP+
8oWRO/rNtarAV1nPACxqT61xLf0qaVG/Fjmms+Qr16vuajYN0DccCVzU8ephZOAK0yfgNOqjXyBc
HskA7ojWNk8XyQGRa2rD37nkDCACCRKaKMSuKrobdf7kr+140SoCCbvkvXKHpGX3uMsDhnqFdlHK
d8y8TMr3WhPY0T9SePsL1uFSUEc+yJ4g5LNBT1c8jzqnnMAG6+SalLYOBXYHE59H3zxLOsB5HuBF
zimnJeOSnQoZowSY4dJY66+u4ZV51m+gkGAlxbLssxDU5vhtfycZbYpwJ2RHRya5WCI8pvX7p0RY
bK09spu29a6RwCOKXUlpOcWkvqtbKWGr/90jqTymkK8rbetzGpXt3R/0tQWTbpPQOCX/BKZOzyMV
isIL9I6NNotLQ7Zr0UL0w1xJjufvuBEoU5W4Ae/0HsCdlNlI6/bUW6IBnS3C6RIR4mratG4nL1sr
jcW8hqtgWdPg//iARMNB4h1beIVMdlrbLUqSLjMVAc+FYzRBXXj/7/xgj421aC+GZKi3GUBUa829
y4vjktHbBFzWEWqOpHZ6kcwU7roohWusZzR4NjxD53asq4+V5coJAe5arxNUwhibd5DLDpHgMtBP
AVdMBc+9xbY9Qx3bLievUUczyDUYarvITzexNH78aE/ud9fhaiBzfCxAy4WR1eqyUZEo6HKhI2Td
589nhxMbkLf+GKadeSyJOT23Vfv3NdhQeiHidVkNUuH84V3BL4Ep8SslGcBlLDMPBNnT+wfjtpsU
1KvlPPZNBRRzXJM93EAkDmDzDaRUwwlJCuACdEZzU+G3vA68yKudtyZ0JudAq3w7C2es9oVpFPKE
o+whDWL89yboXCaNdmCxoRuWaxeyCi7ObLnBLWEfLML8jRRmCXi8dOOe9ETBJdGKpaWtQ7XvNHLy
tL4jgA0l/xkYRWFAwoOgW0OtpVmIKEQ8wufdloXBE7kM6+l6UhGvBUwyNsKIfjUY6UOYL916LfEd
XwlClqXHFwxPJ0xbHTO4+nzArY7BhM6OR29Hb5T1IJcydWwDJ4v04SlvNtx4b8BxkpHAljb5u+yW
qHsRq33yZroQ7huzM8qjCqWL/OgKQxaHBCnvM7bAzRnsmUaLlhr874L04KXa5Y3WrmV+9NMnyIM/
EDx81fZJZ5v83+Z+Lq4KQ6TisiUPFZ/+JSSO2o0EnWSxT7I8A0xt3wgx945qKJ+sv8oGNdL7fLo1
x6AaV0sxjfJWslAw91kE71Bqb236PukDUZeoTsIkWtbxwR8WIziDI9/4e26B5JFb4ChFrddX/t9H
LbJX84xfn9sOX0UZwV9KuUdTY2wk9VSy0YLL91L0zsXtqVkI18BpncCQDTxd5n+FxnvMNtVFEj5d
p0tLNiqQ8GAh80sVHvSlc0aeit0sY+rCCvgwnllauyChjMVcVScN/BIy1MG8HM5uXDVo4sKqLSrr
OlMj9HxtPf7TiEnn/shajcV4CufbYWVl8RVVA+ynfWWcLU9p3MVDwYQRzmNM8iAKqfdsWRkfvrMs
GXw3pYiWcNWfdnOvhuoJjIbX4bPsf9qTffBYBLcZEILsP/GymLkmyLHnmpp52do3R7lctjWXZXI7
w+OMKF2l0vYFJnuXKHrNxvw/VKca7R3D5UW2LypqHBZTVD69g/CZsCbQI5zKfawl/gLbxBNrCfmQ
mXZ6kt1KfyuB8+tto1vFM+de6fymonTlCIHz1/oAPAWHlNBZHr6hVO32Fxjdp5uf6gxFwDAG/Kaq
pOXEGmyomrxy6CEzZ74Bw4IizkClKuryb81TTc1hoqUQdvdZJg9i3YuMNHFCtRJIVZ2H7XV07FHM
G+kE+50fvZO43u3dZANnv0gks2SlBOCXA0pyDB/MVFwZmhc16YRbvLftAZF+AwrQFs+tK+dmlAeZ
ueBdJXFBvfoTnu6qNtjzDaFZxv8s02gYHCGNogh2xXa/5fRgiF+dt9iZXfmgPKC8kZdvYqgv73FG
2QNh7C1UkdhLTSDZM3Acbb9MawB4ljzFWUkBdY0jBAY3QpSBYynnZPJh3yBm4omkEqO6jaxVJNUA
frMEZDH0Td6FimBD0v1bp1A6MFKh3yquo0eVKEeLcgve8ne0Le7v8vSka+k0NRknmVQlVqvaN8cA
EeeTM7L5Kh6ppIyZ5YDts/utk5QLu7dT7B31ZTxhVlfYt/MU4w52fUTu2Go4ILYZUMVFHwiiccYP
hUjYIx9nM0TYrk1DsXRf2MgBA4GwCPyM+RwRFLH0bEogu4xyqQhnmzbZE0XAJJ18bRF9cp9Txmpp
G3fA0GQTRJ3slwPg/BMJvOQ/e0EAQ1MQBdmwQaiGyfY8tqmwny2fYOb3Tns/oTT/LUi4Em+fhTWg
k7/pnZIj7/kjHeVsLjPJZvp7bvFbsqV3X5JopyJ2ddB3g3lGHJvhFUKa/er9SBcXjuedyj/7lyxZ
vHpP3CIdcX5RMyu4wM8KV9ItJwLau8Tz+UiJPSuhkOYH4vqGGoZ1YjQnrqqS287PjatF96w35EHP
aWoZGV8yH8BEd8ezZGZ8q5hZSWaSZlRwi8AlpzMHRq/cY7QCT324kaOL4bIsfZSrkZB6N/LObAir
+ZoHztOao2anQe+kx/X4cM71Ghzk6X8FQKGzu0u8Pb0rf3qbwOttmKmGqEvb7488awd0v1GQm8rr
WgZYKacVl7DeGBl0r5U0zuljZ2acRsnVWCIOvLVBD18ecsOeEIXiB967+NsC46KiieUdCHf+Xk4X
kHWo8vFCEnTjOKYeMeodqkjXWmcgIeu239lOEa9c7Aytz3vTu1Qs8p94aEKjh4+Q3wgv/OOaJ+tQ
TgZp0BiOKtdaU39Tld1goSeskaSJTqX7ExU1W+PUVxPbCvKaxs/q/9t7PhACOuvb6WTHyoHmdILf
gzb0SLvUGMSAM7K9vx2cQKwuKjznPU0NLTE7y9bcqPhwTWNXFwGzQP7Z1tU/BKQ4915XCdVJcADB
NX7ycktEou4itK6G5K8I0QcwE15RPrRq2higKAoPna4g/+XN/Z/I53Fyi8nvZfLRF705T9cKQ4B2
yBhFusNsCoCPgV4QlTlPQ/XvaEgLMygSO4I5sqghNv9AqrifnbvtVh03fobbeQaFzZ6oj82YVUrs
0xT9I1jtWUIh8oDhfWrCdIl8rji/nBBD9EjVnli6cBx1/9GHHOb0ILCOQb5vVBTUKE433hiBhAF/
vRHC13ZaSrGac68XBeFLIlRXQf/qhHruhgDia3kCSZaJ4BUDAC6Qtsx/Jl6+YTIBzIe731E/lfUc
ZPSivPQVOd9ZDggCQqcoxcQ4fYGCmrDMLo8atx9izSB0s0Tobq55qdIJYtN40LPX9z04Cig1nHCj
gCTGx9emrsxsz4BbQMFEohiTfd4JBydP8RslyqY/M39r0e4k2HyAme+IyJEOG7VaLBW4TDRDXs/r
b7fYTVLZkzjZF1ZDIfik5aN34Z38+9/I0mRNN8naYmaLY4PK3w6N9HdiZUVRBgOz5Zs1nSltAbBw
O+u1b5WHgu57kcVlrUy4GWdqO/trrU9y7hqeU2iOpGCRkpeQD6TbCwN6BDg7MJMT9tBRUaQFebk9
nNOa34hxg1dDvXauqnWw3vv32BNCVDUdUmD5w6cJdTrjdjVOFvJckiyc38hoU0qGiWihNhU/1MXE
vipJ//2XpiAwzYNS/x/wpa+eD7s/Z5ON9ki2+EYAqo5qCgesAcmUlkc3dunycm67CRUrcHFVe1tS
0XNAGjcw+OTa/IA7J5Q7w9UD8wD8tbLTkGHyp+w+V+92Jfo+wsgmk7AE97MfIoxVSPdWJMOoVss+
NXX+95Gyqy54hZhnFIZGhyqADhhcFgI17i8Vy3pRYbc3ao5K31gAgKOTS+98iT7406KGERRMYyXy
IdvemhHDwrCyZ1S3yf9SUZgpN0joY3RIFZWlz5+u7YyRG/HJm6On/qumIuhS2k93c1j779EH5BlW
b/toejVk7/jbHTFE7YbyJyeZKM2EjmEOg8w1cpRYAb4E8LpLyK4nBtJkEyXd1isd0YOO+uocRge2
vZrbhfLdXtkb44d4+yRC5rJSFJXD9BtAjPQRfm00ltDM12fDu+q5FBEFzyATO4lNkCmq5QQ9KEw5
/xNPeSGejUSA7EgwG5H32r28EozTxZ0cCOO3XQZEdwJDdxaIS72oIe2vWHXG9ZsZVxkU6CpyXEQz
NhsXS2c1YoZb0ZgAZzLM2M9OtcD4AqYkhLv7gnXPgZLk/3At3zCURkMNN7H5DZRCp5MXwzSXZpxY
0a9NOuQKLJ974btSXExZQQt6c0r53y4haR9+/uodzN8SjJxFyWdLBndKI83RdSHQDyNq08BkwXDN
ofYLnHDu+ahfo7UzFvdxr8iu0gjnZc3zuBJb3WC3VzsogzhTj0qMGI57I+loyD8v6BBpSXLZqXFw
Fl7ve83YaB4qwGSUD6Sb1JnNTwiSiqdAUMzFyHroyhm2iT75w3+9f8VsoHVPyBwzoVYEKJddmDfu
izDNUTjbVzaio6r2U8jkQTJQ1uAk5QUxhpU2HNc+3L3zASSAlocPJDQsz/Tpf10XaBryl6jcMfBo
CrxKrt0fv4Ho8CV9LuTog0tHZ+cjv5lrvD1KXUVjwSKMZYDUbGOxt2VdI1RaDc+fzN1YsH2lOuwK
alyRnEwWS4defakLB00R0dOPGzqRAmCiLbZ98HcKUCUDG3YPpBJe3uLYc22xK9KhEHbvj5u50NpT
+zj66lMj278SlIzMw3owjJdkUY6VsBcPSiPs/xUhV4TYZm7w35rQEA/O+cXscF935pGE0Jwj2QnI
8Z7qvRi8K/7wmbRoEcuFs4EKZDEKOzHl7dTz/qAdD0SvMFZSTyX8G5tWWPhPbm82DgZuRxIBiFZi
l//4f6QXJR6LTBpNuy0J3Fs+SQtM9twl9MzKD/0ASC2lQD4p2OeW93GEqy98au47gYfnrX9UX7LW
osF2wlPBUwG0XwaMYd7MjD59EApCu4PyBAvEp/sUoyWq3GPYfw17PqaQ7guA67uFpn7asImAWZWc
+YpSPrE35IBLoZdUlpo/j6lCeJUyvSOJzUz32Ypp33WxyTRgWUuyaQ+TuhJ72kim4KJu4yPD+XK9
hGENoIw1Efk7ni2c2m6YwKrpm1O1QC8k7Ml9ZGhaSejId4uSaXiHSorHf2h1fTQHVMZsE0FU1ETM
FKmEFGZLfkBTCABX4mgtSV5lGBxtHWFrKL8x1E4Zra9O7WzVHaXXwe2aZt1cXHVWgyB0CjEoMvy4
MYPT/wnbvyoe5pgb7NOEP8vBywGxY42aTlkzb7tcX3pTniDku4CpkgFcG3RThb+ZLs0DJwYaHcfV
rpBNVddMZDzfctTiZU6G6t7cQi4m+cnQ7oo1FFlZ66wtxJBWst8rtlQuxwmRc0qtc4ND+ldElwzE
89sCzllxh0JigxBrhgx1r8tYniQW2ZtcVT08mCNiZ2YWDH/3Gl9VtVXsrbi5PFZx7ehCWij/jf2g
kCVmGjZ1UItedP7Zdq6NiOKF4Fd9UMnKi6A17kjxhKAVYc3exL36b9jbCvHx7Z2KtqQznX9h3wR4
N92rdsw1HAYFAjTaWvJ+4TFYXYpg0WZgg6rkdoLKfg2yVZ74+MWd/FJ1h7sFj0aDj/sdbHhUMPf7
LaW/4zNPdCJwZBbqy+UvhVNIODrKrP/7Orv8vZgiiSLpvIdUA73pvEvG0xl3sX7EioBfC0gQjpRe
MdhdLlNCWV9wX3Oqpgkh2Rdb9LGT/58BPrQlFWk1B8LQtb3bn3zaqYBkc7mq2HKVtJK6kLJ1JFhT
b1DKmqIKo4B6M0bquQm1hT7R31C+sRx4b4AR5IrNh6UdT4/g2W9uT3T5h/A5H0700zRXNqiojutw
57cZbs5Goi78xCqQ1/c+EQOB6lCfdF2Lk2OHY0ERY/Zby2nJd6Y8qHyH8J5QAoqxVgQMolGeWR5V
Pqoje+ywKerYG57YdJ0Htn4Rz8ILhV2hzFdO2NSOdET9uHreTkthzzN/AOSo8JL0csfFmByOGnbM
nByEz5fOcLvX/NxqrKB44l2pnkwhvs/yaXUZK5C+oCH49avKEM/4vMGziZhhdg9C/1q51osRNthD
rCyFetaH3oW/er8Ipsose/AkKx8XQLJglNqhhaJVlE6aRETughmvtFl82q9/1cxbe9W0nt2vELcO
bLQsQ4TxXZnS6kFYxE+F/AmC5CuZ0GcE5f+pPChXJ0Zj/ilKmWpmyeYJp0qIMZ9o7rVZqTUOtz3v
PpsT9+5WfXki/dxVhpkLjoTedgy54b1Rfyv1V147tMWfqlSpRZkyf1lqtxSFfUq1IdgTKGgiNKTp
d/y/pz2B+/DHRRoZraYSZICoFKubTVDdbiSttndp7brfxvywAtgsLvW4pX8IwGVu41tqnOJYzVl+
k/AQ4XwJy+4Z+EAswPar+WmKKQD7GaKOL0itH7SVTUHxitjmoIvZEg+Ors1I/Zhs4ZHRUkkdNS5Y
WVbDSL11ifGcDzWqQAPO9FG6bA0XslPWwVHjr0LkvbyKg0AxdZLb2f99Rb4O92BRkZML/fpgIVUw
2ABekG5LCFK/cFJcR7/XH0A4y/GIFz6TWZtKIXGtvxT42hI/mxZ+8lRbfWmcw1GkDvNulxzJhyd0
HKoo55XpYYwvntcKatgLh97+LnwsmTMfGAs9/tdB7OHyrXxlwsEPnpGkxhzsC9oXB8+autBGV+MY
NDH0zcm7BvWOq52gmGvoQUjOIPmgKKz2K+Us62r2G1K0tR6neR6XXyel8uVZ+wZCgKpFn4bY6rFW
8TCrGxO58cy7OZ3cXjIzfhzBzftAgWCEkBwZ0SuxzSU5hMt6/dBmSR1MMDPwNRXHbnJiQFQZiu3H
Bq8ADLUnbQT4ZUGBiAQgieEQMqHmox3jfqK8JIokhaz2AWkwAOmJQr8whSwHjusBBTB985v6NNhf
b4G9bXvIzIpBzGW36Pu7ru140tFBy6odfxueTpTKssvOzvgDcPiaiBWY2oXlSfy2q461p8hjIrFO
UdsAI/0PTcdj+fp/WwoV9XyTOwOT5iCL08oi44CHrWd/SFxOOgdQRK+l7oRrGL0i/a7QTewtd3pp
I2GEimnbCL7dFZGiQh7IO+8RUqC4lL7hrv0tTgrdk86rt4QiA6Gjh3azB+RS9aXcktktWeXhM8Hh
YYe5tjZAYdoWyh4sgPfu3gkM4dcSZ7drTe0hnTcizxq2J1Zz3wk4JwB9DJkCiFRDi+2P5TmvArK+
uwwPTlR6JFfbzXOxxllADGnPUZdxBgBwwiaHlIfDVU+DTI1Z0TRWJgkGqM/G1+PzZihcflQYguWB
yO3RM45z2rG3D+p99Nti5E/9iS9s04gB2mYMQlWKlRb9tou6IusAvh8vvfPv2EKFRDrXDkjBIl2Q
VepJrXXoaB4Wvx7/TQfjB1ah5fUQShQCHs8eGQISDLdiLvjagvDj/cSvGh7PLL28dTN8n5WVTmwK
owK/PshVLGs4mnkokWmUfv7OUYnRCimYI8UvQlgetE3/dZ/vOA42kPvh8Uwa/1x/8MGMMeOKGEhd
plfoPE7a3LPs2tFIKR1A+iJA3lKGQ9moisC85Kj2qAzpdRxnOt7yG7/kFgEhW1OHWBur+xClII1d
gzzteB2eSBUY0DwUolHRjDb4tMXICp1WiBU/b8YdeaauPPjYtlZW2Kt8HToZ2tFfq8HAK6ORaRs4
/sfg7qX5HDffUXrrF811ZS36UyHCaEbogXM1Mq5M7yVhPSWvVLAnYiQ6sv4s+rif7nEJn7wdadnx
AbZ4ueTxwXr3x4EK/IOasgoexmLrwyIxr6LTfaW0zWUPCHTw7y3apZPr16rDKGi6D9aAgbwR9ZCa
gKsWOcj1Ud6sQbk2JPG4lDWqEDe0CexIUXpuIlpY9qAiJ9RhLs3j9SdnNoF8O5/OBJDrcJ0NtWOh
huQd7ffQp3pTDYp77+PxGjjhTq7fuyJ8Y4Se3T9mDJRyyiix4KewaRFcQ0ZeA1mSEDyQTwhfmcVF
NZWvUM/N/j8/DOXeFW1M2hchCP1Jc2frA4QAvIpE5Ys2/4xelT8xwzuIQHWF35kP1aa+stq0eq9H
qrV8azytFxE8bLkfpJhMfCdBX8JUJ4ESXSm8VjNjs0thTn4l2Ccd4w9XEE01MK19EwwaqMsgM2aD
JfmmQOMiRs1IKRQQ/3WR1RMdDeuHMG9n5PY/2Xd7c+0luP6Wlwl2p3tqR/U6cFCXe9dwh/fHZUco
AJqBmb4Ec7AoAqB9fmqx82cHu7zXOJ0efc0jpGQ+FOu1zPqiBRV8BKr70Nkuj5qH5IR470jY+EpX
asRCPMPnI93DgwwDvyIooGUOLRFQwzvKDtJgE0jSv2bOdvvBMSwR8bmHVMD877F6i9lvKLgx7hBI
In1EceWuv7zbmsG3GxSNKxbRleelt8CfPK3euRnY4rUJDT1wnbMSwGjbNhNEq/WOQNq7ZPYTqj5Q
uETkc/F00MiYDuwcb40fQAZ9ES5L4jCR8WzC2g+a23AH73/L1xFqxtYQel/Zjq0T2OHSPnyFLnGX
MltFPNnhGovqFU+376/F1kV2eIR5ud1P8x7tkepZXx+qdOcWJIiwk+Stu5H+adsOJo6HqLCiJcWP
iA08Jb7meJP2peDPaERUMwWB43UOtnEYdXvuUhX191BtnGKaKaYURG13HmJZrzTyUqX/eqJvQGtl
672r1dy022JApA0twvuYUN/wuzm0wYdMNAUmO1lopp6D11S7PD22dP09wno/cPbKEl7pprpqoaD2
/ZDdE7tcM4NmCCtIMwbewhQ9z7+VQVWxjup9rU6fhsrJU4qMFcOdP3IZ/nmxTQP7645Q9uy4YWmi
qbJxsg1dr9nzqf8DuFJQ9K7rY1JZ3ucJ9+iwAqsIW+GP1o1M9igNaxjwlkSevCQRGT1I4B07+wgT
HQ8KDzGsBErO1b2T7UVpm9JVtsPOfXfJgrKijIDwGM/1xMMMNQi1U2Ve39l9zCj7ZrZo5o5qH2ZP
GKSdITpM6bPT/ZLiRDalu2LkljHiLUigp577EP6ewBbv+TseFso3zXOceB0cF0oQPOSM/m2vPUoe
JmA0L/5ce/Pyi0kPr5D+SoGyiOjGyVgn1wurOtAmLLppJSGNXTYs0kSBwojEKO5oeBV6+fZmuZr+
5Em71WAPEoJ8LJ0Ri8nwopGtjyi3iPqhMDqTo25XrFy05LzQVU7x3UGasIOjn/r0dCGlpvqY39fJ
xVh1PxUnHU+PqJRiB5EyttpcbBiGde8fyae7CF0ty9oOkvGIgyfSzWBubCIO57M/zntEaV7y/oAv
7+B3+rlw63kMuUrYmBUDaSUfEPVKfhqZj2EVREW2Zq6MSBbMRhZIysPU+BPJWAq0qGJR+3mKyYdK
getuAX7voVZxm6IfhLRoHBynZHmDgbHlODmIcmKSayvHY1p802mjevb5X3P6saNFmYrskeb6cNnT
OpEbSq3YpplAP4tCK61h2QFnmf9rWCOPfu3anH3WyEzumooDa6TK/2uBW8f06xqNw6xiuGrqzyy9
NELJKcKqcClev4i+/32DPKwIdUyx6KLN+8cuSPtv4obzF0VXXzUz2WoD5BzEMy/cp1xSg3jkgM4f
yvS695EiHzBMm3abwP466WlyYN1DMiQ+0u2DbC6vRB2Ezxlc6LM1w1NS61JEKpaP6N574YW8wo91
ZWhEmca7BXViyI1QgbcxWD1iFB2fGLpt5yszqxIDq9WF7D7OZYGsqmUF5no1ZTyX9qhdcgMwIt0+
1NnSNVPj8DMAkpkdRpoZkKd+gbentm6Js3HdM2+OfWr7/IqyZdcl//lrue0Dm0mW/Vcq1GFCi1vj
nF0AwUbhjJo9daa8gfCcIg2y27mHf0gOAzlLLziUVKOKf0ytNuXXKBR71QGVw083b4Ak7AUYSjmp
lHy44B9wM7VLgLJNy901AGygxDniinZnKiXzlU7wojq9yU6GouYpgDZAo1e8ouXczXttaRhuZQ6h
V1zuOnnWCeBH82jIhKof8UqExGJOtdWBuxvOuLpi690ziFE85UJNJQqol1iGbqdahXMJ5S7XoAYG
uYsROT332Jz8LlX5EDpFgULuX+yYNYPTneL/6jRAkAosZXWxOPZ9NakAg1w5nnECRzuCerUm91TG
Y5Sp8VS6EocDW0q8FXRBWc4HTGpfI+t8w7i7Z37kUIipq6ZK0zX+dpoQjSGHk9VoQKDopwXrcj67
XsfEF1eb8e3mN58w0XNK9IlmkrVFAcCZ7oV+zSw3eeyEFH79reKFL13LgVxHkj75/hln5axTi6AW
IENzpz4IN4mRoglOEare4Yoco6W0ewJWmVQfzMoJj6alZ6FS4mN588Evi2T8bThF7wQqQQIWKhAD
pFqROiH3joOLmEY/RU/QiVLqhTTlIEwkM9YEgKeMPDMlklaJ92sGWAoiXxRwuj0dZ7KA7bVaLZxi
OOmGCjnhsOxrmgE/UWrfR6cv8DGOhtFIvX2HPUuDtuBDwyVyFcGD6kweItbWG8zYbExYxa2MVTLa
KVrE+3lALIqkiJ8qnRx4v7PuGvp3jIVYCJQdkck+I35SvNcxvzdmEnSyM7uDGEw34VMGhThQ5qZm
p3yUNE52lbIJLosYilumo2d0V8bPZ1hY307ZncyNe3fVgcE1BmvHzkUkR5kHAH1RjzxIlfCKIFfw
0lKszVJ+7oZCqU7oVP2mznkfmA4wA/ct7zsuzvBFr31pi+lghT71UWaWAKUGrSMzNb/Hu1U6dreI
1we3QAvdJqvyFL3Ygatzx+M773lJk6dhWeJrvRdjyeBPu1vSIHY+llXdPUmgpsNeAz0D/eFTVVS/
cLse4+bWCPu0r/g7vng1HuZYTMgCU3dMuGPUkYdKZ5SBim/tG7BM3lIrtquQcO+dimvkQomEmdKm
Pyz52HcItJojTbKEK0wAdKZ0KPNMaOHLywuyhzRpHb5/TQq9ycqrbV8M4Xr/V3zcm4eaNXWcMdTE
hbdS5e8JBNNAXazSmehFVW7sEDMzQTNCO2EBhP+BDPJKg20+LuiQiU+3BdgKPX2YLCLz53FoSpcw
q7V5zuHB9APTp6K0pYkpBD7D+pHnCOVZl5AoHsU7QBchftTE7f78cfYZw5aNRJL687fPGIkyyE7V
Dmd6SPD//HIo/0ITOrHnLZnyV9ebHxVxa3W7nei29q0OVEyDyK9JPA1qhdq3pVNwhKNS/dAg6sK4
W1BFq+ur/b6EVI20cEJx516PBOQG5JXCA3bv6X67p9fsMYpu4XJg1qk0DPwgafstb0s+JORr0WeR
TBTnf1V5Lee/lq6I/vAioKL0eQCKPJA6agNCDY5F2eWtjRnKUPcAfiI1CfHwSuKEt7AmNW4KVeMc
Fw1HohgNU/xkURTZt2urcQk1oCSirbq8UGWwjXQPl6R0QlRtU+P/MsFQFVJmtBMyd2MzFio0Q0bc
RzuKCRNBHwOp26wT4p2Xl/p0jr0OUWRLWcZNfOME3ZaLkNV7+SzJtpuSYhBrwmf9wBBRTLRMEGgZ
BSA/xTh4OHDp1drIeoJ5NgTbJL8Rf4ROiv8t9BI2+AXgRtdC9qDXe9nsLmvbCHYEja1rTZAheeEN
MiRFQElVpK6j/hzWc9tGcswdGysKUa8Uxzplz+njq2s1qszD9MskCFeDsj0OKhfDk7k/csQv1JRW
rlAAdQa6KCs636kk8x3n96JUTetboaI4WyH9W0pPKICIZiHn/RZIzt3AcczABHWpqsPQR0EDQy6C
eWiheqCKvdv9A8wBtgC2NHBqh9Eza/7UJCog/eP/CzUJdrNuxdmUxQBO4cGJFRw0MgIk9sSXGEzt
rsFz1D0Qs+LV1JQ+k5Waq5Dqu5bhn7LyOmhy56BgA2bYJPHduXQg2pnR9Z1+9rn1Jxd5G23TJdy6
hpeU/6OmS1QhWJj9ADjd1yGrVVdIbLPBDF/s7aJbEK5K4r65lcr1t0mX1p7h6F3jFUiqf/3QR9pk
ZSidYEkyx8LQTi5KZPRA2n2zpgFfg63PE0Q76XRzZPyJ27Qy2QRVJ9MKMbgj6sKlMuQIvkpnGH/F
Db8l0HmTha76DoMDzz3AXwwPd0VFwxJCT0qpVpeGBV4heYuYp07C2Yfcq2jfgj4EZY2Vxi/WgmEW
tIhlhJXKAvVKmjAc+T+UABCnMo6r1q6P3+IrVIUmGMNT0DEbObsedHGnj6YlZ39M/oho76HxtfLL
pKMlXzY2FR8XGdBsBqgRd/VwmopsjYMYWy2gJoHxyFxxEzM8HH559Uzi92K006Rl5hyvRJlw1ILf
EjgjtjCjXEA0q6Zc4lXXhYOvzjE5UUcffJizJu8+zjVK4dF5wHHdO4wE3jb3DYlTpDffS7LqNIcZ
tri7N3jACeEJxYJUF/ebWHY4GAT2Kp+XdNLHI0KnVbGhy+qMyD33CTujtBlwjxwJUmEmihL8DVp1
EgUka7EP3ZG/99FcTnpxdWf7g3AY6e4KbibyYu+9o09ZPETAXSk4m+xr3Zzb/fIKhUPnG/duoT2c
2Adti373+XMPI5CVeZGp7ouwt4jSgYIDc0VoAzV+G3cxPJOjgcSxKO491UlZpNn6En/yqxmlMte9
NAaevxexcZ71C25caOVQcThyF7Oaip0KQnVRYYSF0hi87b4A9GaOAbmBZHWtoW4VGCnlVltzc+1Y
qpEreQMjPAJ4qNmN1Yi11PrgbsG+PfdDc5s6nPlxcos4JvDNnGlV7y+3+irDPCwb7wVuK135q1vC
yx5GLQFvQFcZ7wfLN1PykEAF8xZ8beu99dEiC0uxw84qwoe8ep1TExsVqTUAkJQA3njr/z+nMu33
Gk7opGeUUrpNxVm33hqFQraf2rKZ9X//nAmqvYFznbYu1bOObcMlh7/evznMyS9Mxh9a7zXTI5Qf
LRMR3V9fXzSyMFOaPBeQ6OkLGGpgc7GKbPsZlvyEpuEowt9Pg8U4vRRkSYdtiJ14i+fQmiIw60Zh
5UunTqbxZ3djumOVyTmoTVAhPPxE2xT+hDhrzpJqjG+DzeQ7gCr01VyCIc+wB8M4qkL7jEazHajV
PLQhcZ9Y1fYGv2zeElZFCtiV9CtsrvdDkNUQAQHH/EIWd+o8MlVt6E7iMa1Ama7yOxdYmZvubbyQ
s2TBktjtcK9eZySuwUTtTRbVGR58wGVBBOdiszn5it5NwDEHaxemRF8PPD2LMlNPzBR9MYcldcnq
MG6+ABXeoQJ524wMJEULHN9zQ3PnIb52GWp0unv/5tb9vj4jGcDIFf3sQ7IwJ+DCNlK2UkmtSVaX
wDMneOkREmJ5lNWfNIKGIeaG17uvWFZbMlDafyS8rUWP5uOFPdT1q/me1KnRNRrRSh5uncXAR5id
34bkgarVLhojctOKI37WGeSQXhOGmz1NQBqLuvnh5/PkJFZ4Je3tXeInYpNmj2lpJFGUu0q2vUym
IZ1DzB08XQKwQl0koiBoRen5LJ5mgdmbKf7gX4rCbo8Nwfoksf9uVC6Pl0O/TP4oNCbil5p6UShr
+gXVLoWeBgIo83M0l1o5SxRALXmL+HzeyGDxeu6hiR9iorkKEWW0s6yL8gzbhojGAXanQqr+Ez0x
gAN8m7KJ4I/duHRgxTCxHMbz6/DV4SuebBjv2jactWwAj95/r5UjPurqb8abqAv0Ov7Uw7l+e7cs
Q1WDLICMICaas8uF9fe3WUorBKGoOpnSxP4KLiF94ypegO0MevCY6XFGopmJD8q/1EUun/y91bf3
pNAah/oD03mL5wt0ZCo0U80lHJFIS6l5wndF3Qa+bK0M22Eney7paY7j7jzdd6DMqW3o7Ho1G3pX
ypY4ONl7SsG8WNKI4QGrficGYNYHueAgh5Fhuj3EMwsYDvCc4pSi5aCzzdlbyAv6iDmxL1OXG4/g
jVFYzlaWbhP6Jl+sFyJoWkHXkKI2kVQCOQ/7B8q2PP5Bsymnd63FDcK81uOiI9f6qcppp1YNxPak
Qxa6m1FJ3AkVeMGj+hRcDE1NleVJ7+M5ol6gLesJ1DOrfql9DdwlN6tszEDPUXI+pCE0t4PF61u3
V+N/WqM5gILVVFOW1BvGRBkMyCA/Rgo6gMZ3VwxkLMV6PI3lcPwaheuQdvXW5SRtE4wy5EXtUdDf
kJxiaJCmgCxiK/0L9GJ2Ti7HfM9QOTM7IxqpEbqgmtIoxsHXgyHcRwwgNPBaODtZibP2JQPGpy2t
pPMWdPbDNvJCn8OToerHbxmihvcizUPrZbL/cut2xeyAud9HxLDrFjA1n++MSPri+6bAPd068JnK
wHhGMYzoUjOpiIfOHJxxkaYpTsoHKYLbK5S4Wb6zcdueQNFLH5YOa7lSLS6BrL4eADwMi/sPaoyJ
RH13pLGnUQrToOBrBXUR+jqI1/5XvjA7Ki84OIEFPvP+u4MGXssayEK73Yoc+79Y3ls18TDzZEIs
IZBo77H7EWBenkcRnuUMhLRrJ/gWM7vh9/jbN1/PtI1M2gJW84JOjJc52lPL9HNgkG4VsyDxigIV
KDVDKCr0+rYQDl2jQtaB7ROJDCcJkVH9wgd7CKiMQJ9mgFf8DjD1gBZoyRIlD+nQixyGKBgnDLGv
+p3/UbfbnRWx0bT19akbkgg0uBeAkdVNNy9RLDi/1mgy3Cp8FoS3j1p2NxAQKAKLu3QA8F5b6QBZ
vuU47ZCfJIu5018bRkgBYIR+7e0ykh0f4soouvcGghSc4OlEE7i/zjxQcLX4GB5KZ2w/lmyt+VnE
BPjLxfz1o3L30TM0rTKBF+e/GP0C9t7Ibv/ICuzjeCtwF7lM1IetY8LkN3bDI32Kuvzp/lrH05+Y
yXVOM71YJgg3HXOBL5x+42e/EswJVkBI/NcvovHVxiWO5qlCCxBuZspnKas3gSpY/2XiGqfb45gG
yVWBVSaDb36EwjDVLcShth9baJ6WBCdTBnFa/C3jKWa1Nmhz+SdASHO8KxssmCjdVwcrnuofhx+a
kj6FqTR/meWwsCLlqr49zSSB3Fj7IamiL5OhzL0u8QZ7Sv56T5YRcyIQUaj1PhPEyRpoH9A7MH++
KpUA943Tpa/mIQdAz0tm8GKKZxCuJHkPGXcfa/BXas0J8SOgpBd7wZLeZEkgZMELQkqaQFYJuRbW
70ghHQQJN9o/zAvenWC2Hwr+IP3A8kD3Wt2uQkL549jGZ1ALjHuOHGi+wobt6ZYSfBoK0d7T/dzv
UiCXitdxEI/tOjym/DaNLXvr94GvZIAPPX7JUgRziQncH6QW/e6FN4Dg47OZQXuMYu1VTpt0e2dD
g2zIX2Lnjor8DegKMh4IpS6yZiGVDvTwiH4G1zIKhKXQv2GqN8Z5iK3c41Efa6fKOOch4LtDsW1+
biOjYEn8lwct3Jad4ql9yUg5fM+twGoNuRlqiGh0OUJG2JnxyhcuwgOmEtWvXpWpM4CCqnvt8s2h
sxPP4J640aP+hBd3TIVeX16olCPUDwFVPZhgRIFbTM3SjCxLV+FLtBlT1EMwIPwsqnBrOY9bPOk3
TjT/fV5Lt834NDHrTTSTQpk9hJLMXCdPXYEpbMqIMDCY6nc0cKrT3yZQocPKOlP2nvrkQIy99obW
fosGR89Vd3PbC0/D6Wm539JUGBpeNED281iiqugxmriRXcUFaT9NVhN4S2IIuq4Aa+ku+HU5vNIw
StRg1jVgioBxVVRxacvN+PtDxG5zxUYAaa2ADRti+TrxmGeNPgHo01/yhYyNDEMf2unmz0aF5Ljc
VUS7vWuO82cJWVdGnJHnKYo2Z4j0l1KCQXh9FZOtgISoBsuHRAFtctf3DXnhvUtTAWx9YkTx5qpH
CpAoG3OXQfy+ZPWaAtCqDR7JT3xRYUnx6Cyod89x5JQCBncas7IZHTVR3s5aatg90dYn8g7D53ZB
sBx1+3F+PBr4AxlTcoSqAO6S916g2IQneGtL0ZMywktB5vRBTKS0jIiBzxGedg3/lptLFhIQsZvv
2u1ehIkOpDq/hqI+dHqTto2HNleGxcZ1++7hMzP1LL7p5Jwd98osYTYBIlB8XU5esaq96UWmA/wg
TPtwPyE1K3tL+3nup52q7P/RShjQwGbk0IEIEr2LtoerbGliIqH4lCW4NpI1YVijYlRK36YmDvlh
1BEh8ofBNTdznAToBlNjQWjVhYxVcs3UxKYKRjp9Xj7qDhW2Vdux4hhEb/t6jKRKvQvkHD+ane/C
mpDTS4q2467sOZDB6e/NWsKk1aAWcSQxPymcQ6uZR9U8nPXp1gCZ9ln2cCKKNwdw6tRxDiFkh2tA
1aAzCnmUtQPXNOx0IFNErX/8FbiFFt2qIkkcR19/BRc1OfArHCaHgHOLf7FSeBfK34mpokx2K0iu
KMTikmo3I8X9zLNgmjPB87JW7w/L7oJvoLt11TuE1RvH0RAxeIjuePn8Vu3wAJhDp2Bm88Gonyz6
BnzMRxnmnwk2dy6FZJxoHmeQGB4bi4ynA+77iKrasjgWL7WGbeoKRd/GYHwz3xfO3iB5o6b1rtwt
AZfp9WUd8AByBSUZLQHxyzl32xayjF5KdWoPQVdYDChpqaQBF+pJzKbY3HxZqaR0889FnNFJPe9E
ibRzUgMm6mSpdHI36TkKgsUUk94hKHoVpPhK6RKx+nI8P/0g82BZkk66OY6QaCIE8AulDeHXpKDQ
913vZq1pbg66FGzuUIH6GIV3jI1P7IpvgPBU6JKVTKYOEP8igUzUIBMEHGi1PeJNyRRKqG/XCaIL
9kKhQeM5looQFKReG7gajqB4G6HYYxT4TJictiS4E/Ov7Dvs6tJ1NQiP16AOMnky7o521ap259Vv
7O2AqLW33MG3cm3NwIMpP9oSNtmtjJR5iCuaDEnlg6SgnG2IbKaDvFWXF1wdasGIahK5UnIYqocX
73J7BbN1AS8ShQOcwasxfI39LjlTZHeCCVhT4CS0Om2572WSTrg+KmrMPaAz9M8djDnfX4hS1n91
YJDYuhFZjqsaACgs8YTu2CpicEdJtFQUCnXBzysG5PfLxCmc9FB68gcp9ucmHum9iv8QoZ4kmh8y
CgHpvoV1yJikHrGSDIwb8hESbvXRS3pUqkV67ZeAD2HDr4uSpdH7A4YIyaD/KbcMaAeTIPgJZL5I
wyo+3wAxcDJhFWL32R3uu4J7WY02rlQpzmJBDL4FXdI28rk+bRmi5zZ4+q9XJLv50gov5whYftol
reWdBGJrxsMO3DiRUpee3CzvvzfHKMklTehIRV8NHP38a9auxM1/j11wCjRILFt7oVAkBHqwZDFP
SzndHPGzu7TJZt4rNK2NrEXcXcQTGOeTPTPLYbvLXVNJ+/TJRkdPZHl3Nmu51XAv/7v+G0QjLMe5
4g1BX9Zi3/wrL3LnIT11cz1gN8t1Or20OI5EzDfBvRrM1RIy16zC/Z2lloH0SN4BM/a7lyyP6Axt
AYtQNmU3PB83+qv/HyK/fecVT0XYcVpX7pwSu4ge4y6S7rDp2pIFD8F/t14wJ1GRZfAa7jCGxUO9
o6wxeFnI+P3wahyf+FDzig10V0RunqudJ/L3VhFv587JnRnwCRom7E/nZhemoPEUi8lJ86KA/ym6
IXza052tX+hsYj3rLZxi7qzQscekpogBRlgscrtOITUoPZ/s+2OchttCnoGK8gIsnUej64PI/7Qw
45h/adx3ctRnKr4vRE5XuPHRHg+a1XuWjR3JKA==
`protect end_protected
