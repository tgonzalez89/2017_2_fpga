-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
viaRZ1Ue4JfRmlkg9wo8r8xdJZWck06QAck2vAaTj05y48RTt91RBxcEEJPx7w1FwieDWQ7s3jAf
qBm/HNdgNkSI9uR/eah0wnaLJ6UJEKe4zUZFdJCZiewIoAmTcIgkqNcKgmI+etW1ymzVMnx5nUqF
/jE/EcsI5nP81Y3CWDQM0J6q5MCCivHPugI0ycLSo7CVrCi+hsA3zU6v5b+r8rppKI7yNrmtKLO1
LheJ+HnVAo6or9fC963teCcEwGdmIGM9CiBglp6aN3iw9PSaXwgH+ORE9lfK4T10wEQMcjEnFp5f
zf4cek/UmrefcyWy+NT9bciy6fXh3mt8tZma3Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10208)
`protect data_block
P6EwE4ce+6cP2JIDXUqKWMjhtkH0JuXce70JJ0kUiGJPbkTkUmFmiAqbhM8rMI3HHGF/kH71RIk0
QSpi3uYAbMVqA4N5yIZaYQrtFnbNEby6yGSBN5/UGyUR/AvSxUqkb2Cb0++PXl2Lb+/oaxspgWw0
nvV3tJdDSczHxKM5saDk34Wb6sFsk1q6zlmlHVufrqLwENotG3e621HdBtV6dYHYvxwbV4VNeSN6
j1q3vHmGe42Eg9HiP0CRL7MwI5dolA2/F/8GTpnlA0QWG0fMTqMJefHKKJBAbf4wpWRmnn/QkFCW
+j0mpqIzbrNnZftGaeAsz+mUS9TirC4jJBh7CeC8NDRONiBcXcv5ewISE7+Ww1qevR45qtruR5F3
PzRvTK5rOp8/W2For15Dn62YDAj7kf+V7YUZgOKmnTKiCY74U7hMdjVnJtWnLUxjdyQND+frt0Sg
Zo+ybypzRNMY2LExiKayccCLzM2le8/05gjoh0FY53VZ3N7ez2ZgTNtzw9RT0nXOYfb86/R0XYDz
J7V7mF9j/2vgfWrHkG5A0DIyXHBbC1N+3YZjSCo+9Ofs6eF+KHzULy6E5uN6/wtGiEs8a87L81kE
OfHXP67XyR3Z8J57/kOpuY3H/6v6NJX0hYQvWy4yVeEBey0Wle0qthq0R3Cc+j8uCJ1okoe3vzXz
PHAFhYpfuKTFnTnrXLzvLp1lTUHFEBs2lNaarU0AhWmorCgLSdO+kPiSiHMQ3PRYPzTCQaxwOfVF
FSBd8bvRHDZf+/BKQ7/yTTMFNbgWa0HbqClUP3jtjRZSR4BAITXhU0EbC9iOwLmVQz6U1mZqNUqT
vvYencvYUg+p9RHXG76SRTokby0qBrp/bNY2XHEgFmf0nhiUm8bW+sxuZPMsH8qAnbQVmWBO4hM8
lOnLWkRIeWDM02gNvDDMFzmk6T9rnw2bqIN3bmCW9Bh0qNufnjq9DT3M8MXnnDyd5AFwp2OMDdwo
uEJ8PSrTOLv5YimKW5DBjYwLdj1IEsItwHdM5sIiRCzD3QEFil19BjdxPICH3jbzAXn79AlGuCao
1LNWo92mkNMcUCBGQbESVB7WlMJ7ECcoy2pGSPW5Plon1DkYsa86hBtaxH+PcSmsluzELY/fESp5
W9xHpMNW0fL8DiTfpiTqNmJkV1IH7Od3iTdnbq7MOlHmXLKdz+/EUQcQBBwcu77TOmaFhghsW3Be
8anXN4SkgvLz7w/NV8SG1dwYoL4UwWIdOSkQFkbh9nXV1DcA329V5/WBsTXJMGONG5jpZZST2F8f
VV3Y7CFcsQ6J3bxHAthyfMJsy8F2bqqGfoUIgHK+ydL1z9P75K6UokoRIzoxbY/fpAJA7xv1oLvK
J5k0dcdoUHGSF/DQdY+l94gBM8OsPSL4/5G6ONnmLd78soHvd/B/q01dLJOTgY5UfxLNXScNuzVU
ZWGn/vExcSishOrkw9fTayAv/KmBSQCBF0haFWMkg8R2NMu9LR7a8izNh9JJBl9MnzpCF8Io2WM2
7WWcTDIv4SvJbninyiihOyAFxW33PtcbfVVQ6lfFWMWI9SCMzffztLjCzVK5jl6JPx+kTdrQQ+Gl
3BpgoUjvEKIyiwPUilxAvAdxWOjpYLAixMGQzR0ebnK7etUsAS3F4gq0NhuprO1i5yqXprFJCDuB
G+6ypn2JZeh4Yq0rp6Fk4GE4I1LoCLN5BMZgPRIomCB+u0UDcis+7eYuVuUZOWQj2upOlGmSCHC4
Dsg4Fvow8agdm84duLBgV2FqDfLQgx1m9MuZ887TmqntBTJvc4IwCGcbnE8C3sEoQX6d4H34lA77
gqSGdR23qyr1iAAffbkZ9yRelJ4UOUrvnI8ciQqM6eh5lOEavhzuJkzS6ZCrwRsQDCIE3ptMeVr/
sHhwF50D8URK6uDAErOIYSewVm0pXhfb/DRJBa65NOzpxuzcRNAfXoDV4BhzDpjPVcCQLWFj69TY
CmlH2nwv1D19w0NiqOOaxGBS+kJDbuzovTlRQCn6xDFTBfSL+PA+V+Rl2AG8w828Q71eFzyWVxXS
sVvyk1mqZ/t8PgYtwWUPZitjZSZRUMFl4SRvghZGXZuToxuPpfnYH4xmDrGmcBGdg55iG02vPSuf
BgVIrbpmP9hMJBaV8AohHMgLAZBjfHt8d+Uhg75GYfnyBp0F+6nTqAUJRMUNV2vFwPwE6LnGi/F+
2id+eH+NwJDgUmCNxQSeDFWMJnH7JJW6RKUO4jgPEdeu28y2zNAm/vdGq3TuGmd0AYTCrBIZEGFe
R7K1brJa7gjrxWBRm8l8dWZrL7i2J7kIuog9OJnj+HE07bJF2jS/m70NhXJqsZjG1xWD22N3gxWG
LaGrfkNp4hNOehjjxvEaSCM/TO90Wlga+pk6rFeRtxu42OFIula+jkzSNmQ6tH+rju+d1kbTvlVi
Mw7hq7L3sqNlsZOBw2hZoem8gm7GRPRjj7OC42Cyf/nN6i3X3GETzHb6J/Dww/5avDsxjqEF+MKz
nfjJctTgS2i9BKTzXfuLxDhgrM6+Sy4UWaBqIsD8HbCXv98s2cnCKxeok8vXa2Axmwp68cniMsvf
nMIypp9wp2X0wSEeNIoBPRazGGWwnnAwiN4X4WbQ8ORJ9YPZeRfC4D/hrwCCx4EzsYBHjxyw1kSr
bJvest9tAtsSjiH7ImNDifwYadSsg9ALsmGqed87ulcxLSKF0YXx1qgykVGf667Fe8cQQuP+Ic+K
dgr+UZuAH+NkaPqelWIHHie2nS3nZfhPlulxTPMiTquL0ymCo4EuEO3MQw+whCTMq7NuQTaFf2xL
EOprZd6eJiCp2Sbm4XmDtG0WQBY6pHLCZLpUkFBKo/2+xdVmszz/aVy/wlvTp/VqCYl94RNXLPL9
udD5lEpdv3pMusws2e6xQP3WkmpO6XAEBJqnRUxWrjFPNeBpTsmT40/UGx5WJtbPAnGUdqU1Q2ys
UwIpGbeHSuf8qBGtTdbmDMQAO+B2GLGMpwY0Ns9NHeVcytb5mY+wlNTTXMiGnJocbd3MWyC5W2Do
2tTvPbDof/Dt9ZGesI62Si6o/Tc6uABogGDJyQePtu/VMEQqtSVhn2TTs0wFHfnvCSTDZu51Lbq0
mYXIQnu+gQid4PaXT365rYxh5pGelt6I/8r+1qcf1r/YV7aN7gj+M7CphVH+cE2TGG+8mcMGvIba
4s/EiRZh4AuSPnE3soSsW5XHhG0hHBIWmk1CjqhfKD2OH/TSidOpoUXP6BUjBaNngNzFjWp4Ebco
i3+KtL/Rm5YtH0LjSzIpV6JNMhbHNC/1pOqg/w1yCDGukPlRal0Jzz2lMOs7ENx/srk4C4SeZpkg
gwyM9S1elKncj5SFbi4Yq6FE7NI9dMO9n3TeAW3BmnFIi9lBPARcpjUiU6NqP4FrxrOuE4OIOPOp
9hR7bpwJG7KG09/Whq3a8jj+2f9MVpnK5p/hEqIPNfA2uKhIw0N0/3+8pvKEB5fsQW5SqLW8nMJQ
uEAPp+WlRSe/HnQ1b93zwAN35RqYtMxM+yOnbdY3UMisNwDHlnvCXXppl0pbALRZIf1ukfcRpwXL
CqyBWwVAbOoAnBs4jQrZBrGfpZbhMjJH0rwGMtyfvst3SysTTFJyigPBRgr7Yi/DyfKbDumlg6B7
940uhQh0Stbq0vtZzdd1bL529ey1D3unVpI8Taldnu88Ldg7g2aWY1UoKkqV+UVqX0mlnUrj6BBo
yI2a3FRVnIITWOq5vOE1DM1MH02BNZWnHViMQIdFPGKZqAmVDW8SSfjFgtM4tdjOKBtXNAINAIYU
8V9BS5IOmbwrRgy9nJ7bdqtjrHtTui7KMrNa0wSy3xKGp1kLmhqdbX1WDqvO8RsSD8PN2RNqzVZP
WlRMWXNpDr4zdG4Lo+VG8Jcw+8SH2gMRXRDJE4ZzBFzhwBsOELBVcwLjM7zP6j8gVwR1QIFC50TS
9c7RL5uGxHeljq4YWRNadBYysAdex8mAdYAsHntOVLb1HuoVK4xEHv3qB4GmqaPCG+r/JUBcEnQd
vsejbFCa2cSd68+q8S+/7e8DV5QOYdsz/yEQrKqedN2O7i+Y3hw7kSVJK+VQlipFMJxq0PjrBk3K
oj04M+DoIKFmJCTUoGDWbiyvVfU/lrn1/EbfJTh/l0eLHfyksmRiepqFn5m/cFHOhhoXJPsRXIem
Kylz4bhIVT+qFWjbOT0h0D6zSkFvZE8ealvtjzIvUMMt+YYyt28ezRncJ/nIp2Lzc1euecLTwepI
gSSK+FCxrMx2Tr7D6Ousaogz8R6xh3u/S9c9LTemas1BsUPWx5rAvesw12xMIwd179aEZZUfolmm
bPf0DLALMHBl1nPI6emhuN272R1AhfndnnlzqYsbI1IVVNcBAR9AGg/f1eIVHhJWNJH4gBFJ7A5D
dCDaMQO9RP4ajOT86YAAKU4vwWbrsgoKt7nn/1zIZyqQL72bvkbkkodxuyi2Oe1s5Vx4qfEYOiuy
ijN/C0VC1TyjKhPrv0wxgNdtXTaxOpj9h/SEN+MLRXx31ljvAfNbfWa10jkAMy3Em03Mab8aLLvk
I4lLCmMUln0TLk1Sgt0wizwqDKaD0epS4aLTF3aRcFOoH4/Clv/CgXY8WHsiNKzxjPahTa/ns4Md
EA5cp1hf8plrCT+hEtWTdrbo0p06G67hMAxrK1DKKcEpCuUFN+u88dryvYHlsMHQLuVtOTkL8e1L
y1rbOmECgL6wpNnW3tNPOeVGYjK7RFBLh0J0n1bn6RYPsRf6HEVyT5Y12ARgUyh754JFDIZShFa0
2AwGJKmX7RBL4CKA2iFt0cZAfJIhicjb8fVGe4j2XfFR4GkDx0GXMfx1hAeWKsjW4C7IG6QTXxNf
7MA+vGrv+BEcd6EuH6ZnjLNn+8Sx0Jk0x6K65ohRRPAT74auZ2ixikK8zmuNk4zm3rWYmcbK7Don
mEupCU48Fe5wItqHAKkKOY4W5+/YDAo7HlF6u0Jy5BCndG3UGU5iHhOnaZbu2ZpozyW+dcXTPGy+
EWJgjDjELJ5HKj5WyyBxJqoiRwmDI1UAQO6/xoCxNuhAQwTN3dpGHBwJA8897YT8LThO6DepHYlU
OcnrGyz68swu7yCjGjujKRk7RcXLL5+GqtH36wsP3zvQowKF0UHDDRAA4MWGDgOABrVsop1T7B/B
mZRtjalyiTE1NAy7AYso8lRQVul4bvK/2DKAEX4XKvU6HZLMKh1vLJYL4kAXX2fYSilZKkerGWxb
2w5Ozs46zUK4alFd0q0bXrj6NxCeAZvrZoTHjZtVf2JEjZP+UP5LM3QjfqU+K/6xe3JfOQZ6opfC
pgMPviX8zF7qDwfCaohfmz8P321I0kpISHdr4C23qsGEDLb0OG17JVJ7B4Au8agcfOMUYRqswG+I
JhYTvPYGkMxe2HqMi4COD4S8345PiNhKoOmOens5GtyfapWhOCYyY9V11g0b+1+WBM8AbdX0FOQb
UEp+TIcW//SMHfPzSaDCN/ZUMgqBELyndvWPcO/XeJsl5XMsRnXxcgWYpzTAEHuSYwNXbtYBnGuW
OT5bLB8joH/H93h0y109R2rFjjFcJBYO3qAn69u2eqdkUvmJ9pX7bDvZ4+U+kZIiKFo/PjAvwzez
oOlSyjZv/m+D6dK9+1hHkbSDvpZYRM+Wk9Z/QrF2lbD7yH5CE1DRfTMtJUAHEJt+udXfrpu+/dDA
7zbVNkrkm3cytOCUy3TIUcYi7Yq1qKaZbf/i6s0m4tuPCMurCeKk1ZDwNAyYZiJ/pBTtl6xnI01O
lfP1QBrF82StkQuhH6MqQ0OW4PLvVDLzQrsivmFlzca7xsk18rtP7nwUbzQD+cm1ycfM2Y72NJ25
TlMX1pdYat+1qRQBxY3wlNX42givc1Q1BIBSGdA2Bg4aud5SU1YfKkAiSOoFY+5q5gXU7649a9c1
sfsNmZ41IDZb0jZ94PM75JVYQbUt0sO6S/0refINvmyWVsSYpUUv7QbiFnWfO7FzU0RJqOOI5mBg
cSoZtt8DLz/2e5xgJuGnOtVK2DCGJRdn17sBRW2I7U+B3TiCIAqck0dwJsNVc1NaTOxSyKfF8XI8
jW2lH8HQNxToafgtskoCB3uNrjz8UMMKDcM3mlhufEsIFionXaj7OXFOQVbYZ90FEbPyvWYXr9h4
g5rAxtsnKXCjDxXImb1FPvhLvM7k7dAbuwlEHWjGRMesKfD4O/w+flVoMRY7VL6X83eM/4+e2Rsy
1ckhq3U1gtMRTMH2uzg/axH6yeraA7kABLCkYt/DOowrTFy/vQr5pxZ0HTp7CluICO7aLb27hmR0
D/l9wsIJ7t3XiPTBgAqskypolOdAF61afU/NtOBQj3Svzk7sR7n42t61vsR6G2//a67WtRm6mt+j
Fqs2nQ7RuMJo93S9gemdz/HwNRmV4SA23l6KTl3ZTi/lENvwhUd0CDaeozF2dRtzuxzIjyuiX3Ne
azCM/UjcV8cVElDHCznjfc32fvgYB9/+7TOP91WrMhhoQg1y5p9Hl7C47Frt1Edm63vTqdCmEZ0K
n3ReLM7yfXeQAHfta5w2pcajX8HGKi+NYOazBi+fmljg5QyQ9NCgJQOvrp9X1HqvDmy3F9JLrdqi
9yvw76ty2oZ8vQemiMzuj0sZRoQfsJIWiQGXOhyQ2w54kfqdiyqPINMY3I0BL6Io2rOIld9Zw+GP
o0oHC6r5gE7cQEoBxlVgqv/Vy38gG1BtZV6mTvLIBf7+hgI6J9OQRHCL2r5DsGyjsZHkbcWlEsmm
3EB1TfDOnlvBpSpqknwbYIyf6usqHbpYzEu0+C5Po0ucR9nIJJn5eMKf/38CyTHM64+LOuo33l2W
CHOm7sxlebWGMPD9n/2VzIpnMkd0kuJa5CB1xfNUCe1B36fudGTl9CYZNKhZfVcv9kWl4Il5oPF/
on8wHVLT6ZfCCwxstWVHur/2/WvFhbLMJGwWXI9+wZY3RGHwlg7dbLhnGQ7Xe8FsBqO6jvCyT1Hm
WSJzCgiFZTK0Bzasa41IOibNsLqcc14UvFs/4f2M6nVCl0iOUgUtVQSoDG63uiRzj0YLzip4GWTR
nkJ2xyIPQ8Y/K4gPy7OrfyUc569bFPN1m0xM/+hsN19v1i8psQASn/dfUbh9BNiXv7C3jbETmBGn
t9lLDUrgBGosrNXOVVLNBSSgwgpl2gCp71lYxJB3U1/xKiDzOvvdkJMLKKgZW8/fjkHyB9d+9aRH
6Ycz5yk9LYTxDsjGggRiCYk9LRH0WdvfUPkarBJB3Hrh9n+5FULC2HzWZEpYzDmG9Uxo1U08CldI
uV+WHy4galgy5jIcUJIwBkg2VEldhKHNZjcfbVwhrcL2MR3YBTmsh5SpH5VrhsdECYQGRbu1+/FF
h9zv+w6G4diFnySFBBSVXCEa4lOF8SqKgMWCK1pto1PrYe1/02fK1KiOaIdZtz13bqPVY8DkPhgP
D1RrawqUhWwcA9UAxxPWqgagFEhXge/U9LeodISGC+D8+re7dPZn9I+Y4RGZ5O77FvBtcSc7uxln
Rxv+J008c57wcbww3jo4puWsmafAcF6DSTNeKw/I3EYJJBVlREsQMx6U2Q2nHeD/cJMtsMSZenZj
pLrUQJNsdVFOfkU7gBghrI5JctS/DQJnbCHqWzx07/o3r0oj9dPYOWhr8IR5RfkgOgnGCKDl+pmN
fanJRGLTjwNGxkJJIGQ4fCMjWWTN3bN0gpoi9KyzplaNeXUSymZh9n0UTOmkp57UPPxSWEnKM8o6
iNbsIaMHuWFNAuNyb5Ko+t2i48qReM6rnT1UYYs+WqGNkoXEGgSbfRzxZeYzmtBBNXT+jxDJdrGt
ZveKBzbxNh4yFaxGC9BA7cfis2L/eh990HVrf0qRiVI3aYbpfFpQkkCW6tm9FfqFKXZsfC4mUbG+
pyAC0USv6H1Mk64gxSynz9ChYpA92LqRocloL6LBvjKK81C6q4RSlHY28F1AH8fzmrhpW1Rr6jY0
eoDJDHNpXfJiFmH1G6rgAGBvLnUAoWAhoTGMHjbedQBG5U6qE1AshryOM9zLX7Q5GcjOF4an3yCg
1tQhZMxrWIAkuE0vTN3d1dqWum6SuDDcssinhuij6lWYVXcA0tClGkMAzvSx9XugqquBQurLoL9V
AWWJpvdXmWiIyK0NgRrL/eiSAwQwd0IcgtOo4SzsDqgC2nmjvPmXlLHCdhz3ccULwC5Z9mBddo7w
4nWdd8OasdI9POzAsDhqig4mk2LpMSy0XnXDrERvMH6mHqXfXzxVpaoxhyT+BwxFeCh7PR77l68y
aLpzcm0NwRALBXNXHEAG14mbhDZMcrW8+vrwPSiDxFLtv8qlFUL+qzgOC+VHAK2bV1NBssIXAFtP
xykLGwLlulcouSFjoqMyn825KdQzOhh2jT2X2xpXN26cXH4PtEVPHjTfl/zQqw7Twdc2gcEKTkng
puTUKlDFImfPL21FNGT6BMTRrOteIOp7bRn6VA+CQI/VNE9fsLs6v97DowXqum24pRPL0639+LD0
y7/nUBazskh2428DtGWPFwsV33tkdWv+5pgI0FC5oZlhDZ2RHJPzyrLO7k0vc0oqwrBKMj2MotLs
ufLePBQvb7/qNaJSD0QeFT5Eblo46SJBvqfFKd3iQ/sfaSwAB6f/JdHObZk7G0BM5anjMhquq9Rv
KhsDen2LM25C28tEQRMj5qD0kJ3csULkxUQqfKT+M+f8S1WGK+KwQnpeIlkbN9wjmCuN5hHb1En3
JdUm02nL9LXuIDffGCmSTV3cHcsPMnV6NAJ0MaXTx6DjS7+KNWl6vVnoyMTaOdMWhjAr3nwRca10
mR2Obcg1/uhBkFJ2xtuz1a6eEm/vOAEgagR7id9K0MWuwsEk0kfD78hkeDVdJETOyzj9mWH5XMws
SZ6niMlgFhxGuCQZY+7B/84DKM3SUSLuTjYl5mrzuKQuWa14Tpki+euaU8Ri5D8TpSZJMNL1LUCd
DAeBrkJwA5d4B5TSnwzLQzIXOJtjOmqQ+WB+UdALISz/DPD11rANOXkYgpflijF1Ch8lPrcUmy13
/dwf5Qa5Ozv9ERmW3ml6Kg5z3LhNRVlzhOl/5AhXaZ7nyeaKPS5Py0x4eZfkO7nIyLSF5Jbe6ai7
e14ORYPxPrzlOePxZnzmYR6mI1nYBOtWRZ6BQEVPhfH/KoujCCJwsiVFqdcj/CPtBsuR4UOvZ4Yc
03BG2GcpgPTM/g2CeTGJ/nRVVO93WBejTRgAiaeiYWMu3yqS1voSsiRBZboZOwRE9KdTnSfnq21z
YAxyAejBkr9+kfY0VBlm/TvLWYYZvVo1k9dogPgLW5q0078YRQmIXPmMyA1uLOdR2Ql9orRBBmwQ
LBJCDi5ZG3yMdMi5AYkm4WaCMQv8GLePop3N3XpUS2dPgTqd2WRuBMF9W8LEZ1Q5RPkOyAoGJeio
1SNGgLE6y3E5crdr/lJCiLDmbBkfiBmiWDSyi9fG1X9E/KHcGijCbWsJD5yTEwuWL1NfqEMC1hHN
GaPGGuTs3haId+U9IXW3IP3SHzQGTtVE74uHUmyISFDCxcUPRQvvVPLveWFlRKs8MSUKx5lAPCiz
sTEb4t3e4SgNdhy6cZQdypaKSvEPYiHc/Y39q1B624yrIFAPMFsxqDmozbeh3knmkHwBb+Sv1OkO
OprVgAZHu5gyYrhnqw3VBceCodc7kXfL7g88Bt2t40lsqk4AnCHm/6TKs8KNWl0Vvz0zneySjH4B
OfYuCiXgW/9lK3/7vgprT4KUAKREN6HYDyzkvTM1jyN92+3XciNivoKurc28C33rif6Yk/LN4I4o
VKfzjjI7WhSDkoQfV+D51+j40PzfwsLjfO7X4E20426jLJHhA2YJmXz6p+ew2AWT17tW+UvFb7t5
EZxpFXAjWFsJevOcuZVhvB0b4RcMlwbggaNCJ2zv59BnbpFpysitXbVpjr8s9WBACfVoX04S4eEQ
nwJDgCQSGOl1tVRMaAMGTD5ncu4JP1DARohr7cLcV27d3q3oARwr0aJ/qOan95xvMRv7zApj6ke/
wSXd4ZM0ik9i4tas0tMavvcZLozjcend0jvMd8v+J5BieVJNWlN0Bfy1o/rJ48kJ+gQ2SnUHktYs
oCm+0lXYuDnjtjwDEiP5rq3zosPN97mGxQTA6wxP+/dBwjazyVnN6cENq3eKm/uSHjjH5NgoPDRC
fyZj9P6yEz1PLOgOMJ7nH9KSudtwcfRy7TQ/A4zpudcrWrjT+yMoZ78WtprQ6YzwaU9wIc+bVwT5
YqWNOAT+d51PXIyn5exAVH2DgkQ0l0TxT7uXKW+QU4DbU9zT8VsXGkYMLKXGBEPGiUe9IGIE7NtR
M8+AmrYeNrmNtnO/43s5hJgLaB5b4ZTPm7eQIH8i1SNLSYbG0wAyCYjTjZnWUCDBhXU4Xv+X4ai0
emq3uz8N/J3btWEN31ec0wGn4GGAF1XsdUcf4IJcBxXi817ZTUahg6+2PKt3LvTab5PRknC/n8eT
0ZKmcdpjM05IEFry/RVutMb4i7nvVDwCzC0X5OeBM4LJeVeEfaLQax/aS029+HNwbzljbnHzU/HU
PBDvk66cT87TfW1US4BCSReMnFmOP7PE7ucwsuRmFmmzawwy1MGOGqLHh22sq5UUyF6ldHKdHqdT
2+g2eXgujCrZ9UW2Hp7GVW7jeKRdeQ3rfS0P9i28QyI4nZxLO6FAFuRSFrx+dQ4WDZkKfQDkpwlz
I+bzcyvIhKy3Pw0xHGjbBf39oZWiIbxpl7CVZLOwp2uZBhpgFJCbgUXirGysQa8q91GHZs0xblHY
h7cOxzlyboHCeexZfLNXMK+ncckdOwaogtrkGzoWn5mhLgjZcnuomoNlhsLHHdv/q1S0Pt40w5ST
LHXqx8A8Y/lUvtRHBiOEqW/KgBzgO3slcgIEN7spGIT96EFaBMOXyLFSvydQo8pe78mtKGlOAzYz
aXB2iff/lSFBnJ3PQRA1JAjtMa6ZbDVlv7sYbOWribO0r3xSh/iC++ChXskGOGh98jaMcicaD1In
KHNy4tg7NEGP/zjmkquS3pWF/i2eK/zjnfKh83GhQzaCW2wlasLpD8bOhh+6CrCS7EM9ZoD3UZMO
8Jm1VKx7YVRyH9n0NabU6cnhFxedrTNVSEmOCgjS+VfkhOa9I5alqgD6uVAcdkxsRxQQntllhurK
7MQLrToYSAmrxJuuO74oWKNopEIkx/SKw2cdTCfunaluryd3m0XUEboVoSIduUmdgtNnJTqSnmRk
u9jU3MrbQ35nwmKTsTp8lG7xLZq/2uib9i3xVVeIZmpHwk0jQbB+z4fyXiB0tvJ9j3NXEJO6JN71
NfuFBK2BKoQEc4y3RQEVYPnvYjkBCN4u1uf5KM++3aGAkS47SUb36ec6oRUlX1OSIx00c8UAWSx6
aFuXx5EUXTMvHjob3EDARFZJGgAvZtqrIQvxVCWWR0YTWAI2Zn35KqiCW1X5ria2k6V1vY3Pbtj8
Ht8wpYBn56JRE8E0mjaDoaTeyy4GkPmFeSWZGVGc3SmlzlKSf95VTvC5CvoTP8fFOGtfgX/H0E5O
GT4tIzy1pQDMrJtgcMvxFfAx6q6BGZ/pmohidlC3pX8UuXYEebdl/asugu63L8HaL4UOzLL+3qHu
INxHcgHbrb4tvy62bMv2Rd0QiVXcQVlTiZQ8Ohmj/qdmyZiLGkVwDmE6Wv5v8rFBGfXS6I5dIp0H
fg5fP28k3pGTlRhm1Mp993cWmV3SFhf5PVH06KeKTa4gxvM1C/C/Qj/Ttsn4+kwUDlE4T+uga3m2
n0LNulfBQgBExrq2+T4Vgdv0Bp7o2WswqxM3esj4z4xcEdIe7uNFMMZ/0b0kOFEcBdb5MWO0ESU5
Rk10GCYaRWHKMYBGNusI4tGYzwEZLPwUivgas5z5tKN2vgnGzMJDeehORsTfTzgsWNUpRlsNKBLW
bzSZI9ZVAZNBPF5St2EQH+uhGxAWq5tUtFQuJZWWbR7EDcUir7xUumlWlloy8AYgGyAYI2kxDh+X
Lecu2KMPu+psaIn135AWDF6Ep2B4/Y06Uxc/tYxxn46XcVYIXyx/G0Wob40G46VMGKU39Lo/O7Nm
mbK+Srt23pNiZ2FTGM9Hi4BfW4ywFO7jKNecMCOqIdxEWjPDi25EGdsGGpSwqKLEShMnKtcJOkMF
YdxEr6qZUmHls8umNjVe+SsK/EB+AE9n84aaqOemM+w0/PqFtOTOHoYhQcNK5nfEVeL84hgEgjPl
DNfNUDaoTmGo8JV1HgGGnzd1ekHm0z9ncXuz+32YTFd7sjEczT2sfYfw7qUXpUu82ui4qoEnhZxk
sKLX4aPFeHawVBM8HS3btof/8ah/VYtsRRvxCrUDxUN+GTh+WW3aSXbZFIyJQEKRb9kdTDqD1XSs
hagI/LnWPap5aJzuM+6ekqoal17Afz5/OGLrwuK2mvdP67O5aNT/feb86kBUgPpxdzcCtEkxwl0m
WwVcK9tfTtZcpwg7YbwOrlga6lnerWCR5vlx8l4q74ClX/dr5Mgy0OvVHG1FFNOfo+JoZ3166LB/
R2ibdPvFUU6LhVoJCX9qjiew2V/ai61DfVoBCpX6lFRq97CeM8D6tEzcDQAe7zhuuJmp9WuE3i+2
bTDfMwBnPeV9p8msDEdbij1ZO2P6gvZVbg6MHx2AoQe2w90yuHC+rrHC/aBwvL2h6uIrFjG3HgTG
nTJiGDqtxe4zCP17HlayNHBzsPVo8VJBOpiY4nEYY2G5+wSHfiZi2GSJmd6dJ7v6MZGCOSrc2Zf9
kXg6O1VBCMXmdAK4qNoNg4c8455AKMENBmUe2Iv9cSqPxlNt9ZAXl7FVnOdAOV6Jmo/bi20fVc9N
826Gap4B5H/84P2B32AUv7CovbiGKJCkJoZLb0AqKYbi92Mqqb5HwxMW7wBi0ZidSYTAIF70vRCm
uqvwazQw4RzcJ/YKCbHkMyXzXAqAjdFC6VXzSf+rDUpNYg/HfEo574U2gqFNje5IDp/lWgVVyZ+K
psZuOAXZ5P6bQuhBVTEAShbujAwq+4ZnKBgA2cQ9oD95P8k+dNdDC3E5ei6bijSCsRSnmywYQ1tI
TBGEvY0Yl0dabtqbhi9CkJmMi5a3zXW0MnQh9XfzjrsmC2TOlXDwQxJpbJdFz0pw0sK5vKALIdaG
6u+FEwMm837Z6qNSFhvxSkCuT41MpHHUvGMB5bA28xKgB2boKrMmk+8W6ATMqRjQHoIxrVt0od66
NANG7gIgcSnmr4j61226Cd7cbRPELcfuX80uNYaD4l/Bj64DPK7RCpGyH2/d2cD9Kmr/1Wduyqmv
4yuwGRrzamaHyHRrb9++oEUDYCTrQAATDEGV9cz0UhGuRtcRyX8cLjRzwfv/kZMK5EEba/bGeUVc
ee1nM/qBab2EswsbYsKcnse7W0Ay7x9xg71CYcot3xIAjEK+rwxXVFV139eQVlw+ofuRmeBB0Yaw
AUfpJX1NWmnpZkU/JcymypQ7wUcJL0o1+xXP48XIGthuHPC7OR61C6G4bVBtHj7xGQcHTq30jtXW
GQKV64BE6bQCuU7O0D3diGBqd/Pjhqz4dnaNxtG+kDlaXqtigCT9NBFX6Bm4ohgltRQbRNppawvM
4VVfeAY=
`protect end_protected
