��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR���[{�T���CK��TC,���:�
&��d!��]9�'D`�"9 S%�aQ�`!�6������V�W�l�a锦E(�\gC�slu�4U5=1�N�m��l�9ў��P���B�@+yg��=�}|֦���ָJ%K4+�����Yf;Y�^M�С�c��ݽk߇���[�����&�4��,�~�����*!���q�6�����w0ՁV#���$ݹ<���}���w���}�z��XҒ0����f?	&Qز,	�`_���E����3��:�/J\�a�b���H��=��z9EV��!4��ح��d%8��]>��'�њ:ӚzV@�4X�SX}�]�fr����
����`7��?�ƾ_*���یA��N��Խ�|�x��d�/C}��'?��˘~��;J�ܘW�kԿ	Q#4c�\Z�C���v�ݺ���4�p����@Jb ռ�X��q�T�9f��T�M�c�8����:����Q#W �uQ�:��7��V�[�H�҅4?Wls��>��4`0Շ�y�����
���w�(v㓯0�Ju>[���v�@��}�F��%�]z������c�f�TkD,�~8�A���*��$���u>�[<+P���x�Y�Y�	��3X"��&�Y��������L~���bj�+)�Jַδti�:������1�*s#�yO�t��7������~P,��Q��6��1dmi��N�Fe��kz	�p�T)O��v)<���ʠ3�ϒ%�H&�MZ��������<��U�O��r�%����)�0k����'z_��#��a%z�X�9%���)r��/R�� �hH\�?Ix�RPpW��]��%7�
/.&�H��(j�u�<�C��p���n�նdAf��.c[�ڰt��	gT����D�Dc(r��}Y�L�r��e0C&��U���)T�=���{�@c����Î!�vY�%��n�ԫ��M�w�4Z*�u�;0�=�8�U�_���;2��do���5�������7��M�f��k�:H���&��u������Á#�s8U������u_Ҏ�ڰ/\�#PD�O��o{��R^9��?�����������^2�AaU6���i��_@\�6�n�j��V>�m4��uģC�_;W�1�ŏHU�z�d��Fʢ�Kp~�q�aC���S��T�@Z�U�vdxX�����Y6���m�oj~o�O��u5[�����������X�����}��G�F�7���|��*��ۉuz*��q.�2���er��`z�w#�~���\��*�C��`jD�r8�`��G��W�v��d4:���e�*W�Ԕ�wc3��a4���Cz{�/��f��H/>o�H��_�f��8�1�����[�a�3<��6�G�����J����w���(=��V��Ѹ�F���٠Y�K
39��Es�#
^���Hϳ>�Y�w�W!h~~/����M�b��6���N����  �� �k�o:5�lBn}2�v����۫CFZSLp�8���k}��l�����K���)��� �IK�=u���(����c,R��uUT&�WO�VA�����[�0Oã�?A;U��������\�8Rz���2���z���Ӂ�(Ed&�rpY�M� |Ž�g�di�'�;3o�cc�x⁳�-��Ux!�п7��i�L5y=��)��z'���Q�"���]( �t^q+��8�T��k��]*�0^I��I0ڝ�0�"��
��
!�
D�=f �E��#��4x�1>�:@�VU�I��CwO���s\�:i��j��zX�������XD��P�&g�k�@���:�۱z��!� ��ˤ�sY}�m�A��OO|J��`I�+��/�3����b���>I%<����C�=z%EaהfV@����?yn�Z��U�v8bM���3~:ne�2�ǈ�]��3HL!Iu�y�5N�	ǀ\�J6���6�(eH�b����S�~qg:4������w�`{m����o���$R�Qw2�[_X�j�[�4 ҏ�/���Q�?�	�/eб���QH�(v8���t+&Çs�m�u�fs̷����e蛐f�H��:x� ��oܦ�VhUoΠ#eQ�����/��m��u�����3e��v�
;��D�l=�vf�&�U���W���uF>�o4n��W'����S|N`��VDvb���=.�I
{���ހvۜ��=s[�I�b��1X2�J��?��.uTJ�3�Wo>:�����(�Ҍ��Hk�X9�҇�K�8�� R��uq����B,~,��eُ�>{M��}El�߄�~��K�jH���5��2�[㒓�\D�h�ÖM��
d����'8G"��́qǅ��+�t+Og��;>��m~��E\�c �q@1�[�b�HR�\	Ϛ�ݕ9�S5��o���w��F���fg\�Ԃ��/�[K-l{UP�db�H�/�^��܄��^%���~J)��������e�=sJjr�,��"�00�O� �U6�x�Xƌ%�\���JoόV|)����`�Z{��֜��2h��ը�Ε'�MLaC��Y7#�
��j�I�a��Q1Ǖ^����D%U;����>��磎���)G�y���(��s�Dת32�`X��2�,���ju��#Y��	R|fp`'�\r�d$��S�3�32P�˿��!睢�u,ji��Z�3����r)����T�����ؿ6��i�f1�@(s����6�R�N����P�N>E��X3
�r��������߳�^�̺��y˴.M�e�{�>ym�]_�y^��k�d�e5���,�{#�Cf����ns����b��nӕ����q0�7`�R.���u�{�]����ڋ6,�������tV�M)��XzV�1"}`�c��"��B�C�����x$� ��:{N�*m�AU��*�U��>v���8����V����lB�?
����M���/*�~�]d�d޸<�69@�a��=�V]�KF:Lc�s�f��1KE����b6�$�N	�}!���9ˣ
{��ߴ�|����ijP�G�ل���H���*������i��W^5`�eg/�.a���yDa���=��	��
�%���-� 6�̌.q���H��nX���A��ȿ��F���F�m�Po<u���`u��N̴����%  e�]&5ϳ晪�u!ĕ��Op�"�!�\ �[��^�MJ����$<:�)�eK�����E�V>�l=�+ko���բ��a153��d��v���"nN�yT226��) ��De/��N������I�1sTN���!E�{��_t!W[�x�ҋ�Щ��./ѱ{`;S#I8��z��w�!9ݏf�s4��VJ�a��4Q��h�����<�T�������
ǳ<���O����=n����x�&�c]�t�����>F��@���@A�12o������+x����(W��!�`ŊLN!�#���^�6��Gc�[��?y�����m��*s���|����*�3��`oB�?�J�:�fAb`�+F��C��O�O
>�RTE��CA 9�֯�L5_>cNR���&׀+6�;[�Unp�%�^��[��@ހy&o=�έ���к�����,�s��E	oӮ�iw�g�M���P)zS_�a"�s[��������"h����P'�)Y?spڮ
F_y\R�A�� �`h0]����Jt�q@�����'J��������,gA7�e&i1Wz}i�CG���85m<w�5��� Vw��}qp�i�Xbһ�)NBϑ��
�uJ�$�L��o#��E�,�9j��"S��b,��}-�Þ;�T+bM��`�oѣ	�����CZ��)]����t��t�� �<�l���3**���˰�$�ӃԵm�Y���L������pa$Y%5Z�3�l�[��*4���A���")x�b�g�6���������o��=+=�%�ҁi�Љ�O��c[s�9b��8um�4�S�n��lRCC�1T��z>�o�u��T!D\��]Ұ�@�*�5r�|G ����ؓ>!F:�@�S���Q�`���J`�� �`�Q��E����X7��eyg9�5-��O�����,��hTx�ty=�k�2�R&��k�7�����x�xȬ�����T���^�oO;5Ei$���{A��}ƙ-M�j<�S��|����s�8t��l��}i��Lv���E��cHA���̽qV:l5�����$��8|���Y�=���Q���_Ԅ�D�C$/-:�,�Ĝ�5Lz�(>uK�ώ}��a��H������Gg-����ޟzUva��X���1�}�(��<���eG�gV��[��N8x
>�ר��2l솂7T���N#��rp���o;S�g�x���~[cO:uLA�,�#C����S=F2�{~�&O�t��F��=8Qs|{n&�CXC�@2�>i���Euxp�­��!�qP�2x:,�&�;��md�`����p�˸�ݒP���5�߸� ��7 |fW��jNh�;�h�4���O�R�U�ܲ+�p�^�h�px#���)�����/{�U��Idjɽ
��t���	�}��U��=_��헷*��A��}j$�	nvY��"��C
�0�|�m| �!���,�8Òs�þʸ��W��=�����İ#��d�BTu�^^� �\)o�(��­�����R�����X	i���ҿ��mP�sE��PFжe��u50�B�y�m�c��U�m�~�L*t��d�������hh�rf8���;�&�f0dak�
��1�4�����@kZ��)w"j
�ڡ����7���BF�n��,v�~�m: �Z��J:Q8i�Ҋg��G��idJ�)_B*\�`*����E�C����L�e�VK�� �[5�ݔU/ƀ���0���м~�W0�8 �ò	S�P�=j�����X���׃|����R��ή��@�a�m���.�[��u�G�`��O�img�(P
�v�XfG�X0ȝ��1E�������8����	8逃�y�њ��-�;�^��Pc]��>/jvgς5��Ć@	���{��4C�j�TwG�ݗ��r�X��uh@�1����`��&\��EXR�ʸ� ���6�u�4��W��D��_�p��~J)@����>]�`(��9�1Š�}���W�F�~����\���($ٹg��m;��
�}q��N/���e���o���"�z-R�t�8�Z�D���M ��-ז=+L���	2T��:����:U�I�Zkv7���h��c������'E�f��,*?9�~R�J��,YV�rn7�2��5Lw
��#�QԮ��)�5���&�8��u��׈��F�V���ıA�+� ��Ee90a*��z��L��8�������{	nq��0�|\<���ˣ�_1Z�w�<L�nk[}/�[\������(��f�$Af�2��SI��1;x�1��|�ʔ���Ls�(O�`i��?��AS�Jvb��#���j�)/�}N��o��a�Y8����l88�ިt�^u(M�G&�E���VU嚭.�cy�cp�Y7� oW�H)H�h�Gȭe?�E�+2��`w6&j���E
W�+q�4��",^������"Í�ƚMn��F�e��^<hMb�vR��%�R_��/#��'�,�feӗ1R��G��e8�&j�)������3�J@t�������X�ح\����(�� ��ޜpJ�k��$V�'08;��e�U�X����uu�H<R��ع�X�V�_ׇ��ZcַI�PY�]�n��v�����7�s$<p�g�I,"Bt�%�;�H���o�?���V�?�|2���\�F�p�M<�&�X>��rQ�D�S������.���6�Qv�#:H�X��P?���m��^3Բ��WV�m��R��ߎ&�"h�&J�V��U�f�'�>��!�2����j�8�'z�`����Q�"��K /X�[�ux��/� �4���w����8��yh<�+��
���V�-��|qb��(s�{�6[����U��ʾm���%4liF�?�ib�͡�6���&"���r���������d��0\�]��ȫ׍��ԙ2����%n
��F����70�N�$�E�����y�����^'}-*���E
�C�|�Pd]X*~r��w0�E��8n�E�ǽB���$��0����;�a�&�#Atlc/��ZS�k��Z/WX����W�}v�����r��/�ĉ4�ԡ,A0��B-3���,ڢ� �t�E��B�,m2G.T�7�ǆr+Z�z�DJ�+��a�Ҵ���B�y��E+�՜��_Y�lj��o�2���~�s_���:�۟�\D#�(L$S����.�h�n��(= a6��!wz��y���� W����nZ������Y�PN@��3ߍ�i;�:�d�oo]��`z+�
1�meJ�9����e	nd䝯*����`�¤�]�e�;�iX��vy���w�/�y�)�G�r����fT�@�&��I� ���y����������2_{�r�g/%c��c�����8A��g���h�Ü�$w���d�r��[��70����.(��Gc����)��x<YPu#x�@�Y���1�~�p���񺼇L�!B����x��-'����U9�<F����B�U��N>Ώ�ڧ�'\]jl�o�r�IU�k\Y�R�2�Ox2�Cf�3W�/ѱ(o	 �ω��-UK�8��Ŕ�&t����[�Q����;;˞=+�4�!%&�E����tWᠶ� oq�Z|���Q���.(~�U��g���µgc�F(��Zl�#$R �B��d%JC�$S�b�܆�h�T����0F	��Gۺ��=��������n�Q����H�杕��Q��)��*t��}V!/��	�?�@{�B���h�
r�G�X�8}�yŊD(@�$h��>�$�D>�f]���D���q����\��k{ �Z�aiut�Ͼސ�ȿ���U�?R��E,�?Ûu!@�����*T���azWG>�wۜs��������$4TQ�Sa-1��$��:e&Ѧɛ�NX�YO�)_��P�b��Ϊ�}�+�ȗ�);�Ƙ�J,�XKV1���v��>�C莛�~�|��(�HSc���Tm)�����|�j�,��u��Y��|�<��jUz�nՔ�PIj|ۛz��8�d]�^ۍFdX�|�#N/�>,.�/��$�@혾����<P��&����3
R�`<nph�l��;Kc����M����hu~��7H>"�(�-]�P��"b�~{d��0�B-X]�vy����\�B�Z��WZ��O��v���i������t��WW�7��@��dx	����<~�K�?�a�Py�GGq������=�+���Y[��'4�+0���5�S�c+��NԄ
$.HQ�v�W��-s5Ya<_$�1�оH�u84�C���;������e/����N���S����e�F�� ��/I��8�s!�$Q�M@�Ohf@>s��W��u�*V����/&��u����#�rT��Q(��nP�I�C�O*�^�J��F�FO�����X����!BP�e��m�@��Ӈ���Et��P4e���W.e;�i�Kl3$hU����J�T*���S~*���g2�{A�Wf��Yye�^nJ�+B�c�^	��>:Mx�̖�M��_}xK7������K!�j]�z$��X���"o4�	�� �X�f�K�kZF�f�a��:���,r`�6 ��нX�~�EE�+pϒh)�TQ�܏�Y�4��60�@���Bo�ʄI����1#"���54A\����2�e&�QM������Z�E��u��}���S��\Y&��K��v*�a�n���^���#m�~��S���s�}H�ell��������|�XZ��{��-�~���̝#�dϝrS^���[��%a�p�%Q��u��7�
��$ �^3���\ĺ�C)RS<� 8F[����0�4D@M�/D�`�
����)y�~�75�B�}��3�H��F�i�*��}�N��z�<�å�	��u3�7�t�y���u����U$d�X�w����!���S�W:���P2ħ��!���$xF.h�����	Ԟ��W>�]�������;��I6۝
�n��&��m�@шk�.�C��θԬR�Y�uĝڤڈ���CU[��~��`���D���$sd[W�Q�']�L_��K>�K.�^�E$������k�;���̥uZ0��Z�s�	Gكy$[؈S��Y˲�>���5�3�[7���~8)5�mY\%�K�R�~�VCױ�j7�&W��+�4l,��#���:!1A�}9��	�o��QwX=���e�FF��9�}�!ݭe��'�V����b���N�OگW��t��v����Ï�V }����㋌.bZFՈ��yD�H���+�/f��Os9�+��YoS��uy}�<Rkx�����b� ��a hv��u���ӡ��Ms��Iz�f��I�V^��5J�'�7�|�dJΨC㎖7��I��4�`a��d<���ȆxݧZ�:$	��1)Dv���՜�}�D-�� p�,S��e���.Q����coU�0{����S�~=���$�$>i?��V'Q!�D�O��FOE#�y(���O�O��J�2Zo"F\�������"t���$�����茈e/y��ᕪ/�Ϝ��a��2�ڱ}~1�eI�����#������e#��Ⱦ��bF[��uL]?�ϵ`�Y�0��>�o	���g觌�`�N��n��g��)���]�P�ʟK�2|�Qj1���,��b���r�\^-��VM������tkZ�޷�-L9��h�j�/�A_E�G^uNkœ��<�1%�ڴ�bs�3�VN�[�mj�e�x#j��AOiFQtdp��9����*�/����:?��7[E������p��wJJ�C�t�~6#�L d{<4�"nj��s.x�&�A��%�Y�	t�= �>VB�`��i���19�l��1������F���rJ�Jm	`��~���+3j��+#��n���u���Z������Y��3�<d!���2��)�ڐ�1S������`�Ep���u��VBwu��np����3Ǝc�|!0R�|�j��W�dA�fvz�܁��^y��T�׶#3���=V�HbTů���l��Z����X���.l�bB簰A����� ���3f	�"ϛ�� ��ϥ�J5�.|��;r�)$������o1���o&'�Z:����Q�@�.�,UG<\�ڌ)(�~���t��w��/����a&_�]?�E\"�X�O�F�KbF�᥋�Q�a��&�u7�¶�н�-���R��TƉ�Oo��ܘ���;�q\����P��@���8a��&YR7d������a��f�� K�'*������)sZ���$5P���R��_������k�?UrV���#�3_�-�h�Q��0HTh	`��!;�ÚJ�yy�Y�����U����zK��� X�3Ĳ�I=iJ� �Ȫ�O�	'�~<y�lJslX�NIN�g��^���� r��| S�� �GOX�(>o7�^`v����2�|���i�1-iu*ǫ��W*��oa���Q���d�����s:{�A�e�&R�^v#]����xy����=}���6�,�x`���;F����8%;��x#�6���	�J_�o���r2z���4�8�������)���_f�2��׬=6���QA�S�J3Z� WW��0uP�߈�}�����,�b�/9J#O,	�%�$��ۦ}7"��=�����vӽ�ON�*��->�n*����Ed�%��R`� ˞�I��^!�~�n/�#֮i�S�9�=[?1�1���+�P\ԏ�s��l�-nV��.)p�(�c����᤟��ԅ��9���~k��A���!��l�=Vcw�-IئSޗQG�w~"�������+���TW�A�|h�J^�0�m𲅗����(M�18���M�ŀ�ܩ�{'�+�U�_�����^��{X�I��%�f��i����� ]��<:p�´����An�5�~a���m��J?i�(��"֪��!�^.���H���� ](I��:�/-1?	�-��.�r&�j��U�O��,�Vt�� �#�ep0S��*�ye��JY�6?y�ᚊ$�ɴ?hݯ�����N�P�{x���|�3$���S�9���IS��G�}�k�@O�DYg�A������j����Fi}}���o��w��~�i�R#%}�I���G�pbcZ6� q=���!!����Acv������t:p
~(���8�(�
���Q�U
�qȋ�ęv�A)��4�`2����y�w�I+,�T8�ſ��~���+Y9C���*f-v�Am���Jh�"�6;���'�l��V���W��ķI�uݗ8G�ȯ���"�BF�?��'u(9�
MZ����03���>B4A����e��k�xF���Κ�9s.�j����۞�K&{3�wX%$9N���A1��e��f��<��}|Nrl�QYC�:�#��Yf��ȦM��p���5�UL�0��1й��9����fb�9�������aZ^�8�INX�� A۪��-�yN)�+C�EP�C�颍bH$i��]��:[��kHSV�Y��v^���i���#��oB��[�G�#4d�pK;am%�vm_;4��w]y2y���(���k����W���$P��bj��H�u��O%��;S��`�sU���GX����2>=D�=���lT�����rG\���c�8��z����l��;��+�=��v\�ټv�N�Q��K�_r�w>:��M�
#����	�� ���\M٬js�p���~F�.U��}��O��_W��'���<z� �۠w���ӽ����VER�^��(`"������������ ��r(r���xֿ/��}jw�AڥQ�;�#i����y.�6�����?,9�T1���^����v��x�hY��
A)�YV����H�#���a`�wnk�B�j̠pȿ-���r�0>�#1��Y��,���Kک�(�_S�OrU����bbr��L�w�2HT�3m� �:�'t�}��m�#��eK�=`�T]��<k6���p�9�h_08��|���W�-3�5�7(��]T>U��&ʁ�*�;��L� ��xa&P�a��:7tC�	p�#�I�&,�$u(BԻ���y|Y����6W�����h���5����-�#����`��!kɴ�=t#�1�l��E\��g|�:B�6�� k��%09�m�P�Qf]�E֔a����s�t�Uː��(��A,��X�&<�.F�#���ѫ�H�T$�6Qc��#Nu�Ě�(-͈B�OPf�1X�F���z���y�*�ԑL��5����r>LM�����F��8L��y*�Cu�Y� �6� |5l/�S�δ�"�9�A��G�Rnp��h� CA�Ȍl�2b���2�J��퐴��ET��G
94#�ͤ��[������������֭�'�2a�]���.`�t���;·�^�FK�L�����X���l�$�{r��&r����X��Q�8ANl/ם�xT�nu~l�x�7�n`��3�ľ}��s�������ָ�������^����������U+Q��J@��8d3{m"��R�aF����p�:w���x�T�M���� �(i�%�_��U">]z�⧪:+:���M�\cO~��dd��K~n��\5"<�q��w��(�ĵ�t-�J�Sg�Ml�c
���ܿ���l��M�v�k���2�H�O��k��,+�����횫�{�� %9���+�M4���M&'b�m��7A����~d��f�֐����s"z��M~��j4x[�m��Q� �EP~�6�k+&C�+4��PEɿ�<���+�1̜���%��m����淨��=�e�,#(����>�6IƱ�y<#�*JF�G�-Xc�׺C�o/ۣP|�����8L'c��(����,�Hr��{>�nU�Sr���"�(V��ަ��3�%b�˒�7�*�q��>��'߻Ql�`�$L��ɱ��o�eԾ������9l����ZPJuơ��r1�#��E���jd���;� ~�>Od�$�yr���ڕ7F�(ZW�Un�n��9�&�(����5X��Y������E����fa	���\��W��[F��u=.Vw{�;F��":��9��*���f�j�t[�pp�-���q>)69�mN�Ht�}��Y(�˴�QK�ݕ|� 0]�À
0�a�������o4���,�/sw,��e�D�e1
���ލ0��������8F��wx�D�98"v�X��̚�=�d6&�����fUEK�ۃ��>�^���N2YgCxP�U��`�H�P�E�4B7���f�%����'�k/�f>��@Z}�
=�f�"���p[�!q�����k�\�8�e��gcg%��YW��]9�|tT��O�#>.^	��%s^���)bQC%�����K��x�|J���Bґ^�������i���s����t�.�tХެ���`⤨�湰?��N��<B�<� +��so��8���L���Q��(�M1}��]�Xa:��-p�W�2w���0E�s� �n|�Gڕ%�1r��+�ᑊ���Ky�RWm�S�߱U�D��6��潞�sc'�?wS�wzr�8�T�&Ik /�}�mi�v�z�{?1�N��k�,c$,�´n�4je�L8�j�ۺ�(;GE����e�����<�b`��
�l���7��C���p	��E��/�� *�H�^:�#��^�~#�셰J�ff���q�����"��MY��u^,���ē3��N귆A���ݱj6^`MFA_ʹ7������b-�)`�#<ŧA��T��q�C�[�2Q���6�>DU�_������Is�^�T���:}�g�n������ �0T��=�'^�Nxs�ÐBg�{�E�*�#h0��M�$�Q5�?z�b��<"[!��ؐ��f�$�b��MK���%螫 A,��KI���ϑ�0;�g҆�"���RH��Z�k�ږ��k����V;�+s�s���P��Q�{z��!�Y�&��l��,|ʷL]p5mj!#�yK�L~��n1���m)�9
���+/�z�u�������I^���4^�ڀ5l��0E��7tE�c͓iS��fD��'�:X˄ �T��<��;Kyr�o~�L5p��.���/Q�|�@*�b]#|����>͘/�x�4%�R��qx[�@sEAQ,����2@�t�e�Dҫ֦*s_���8�ԤnɯFݱ��4)#9fpi�5C�5̟��u�9�Ud�e~����%a�+���F=`�كz�]&�����l�8~q����vM� ��#�q����=F�tB"�Ֆ���3���n�]�]�6�npI���v�H���r��L����s-�m�����R�,�d�P׬�6-{�}s&�	G����<ۤ|��~�?���S"r�_r���O��k�n��Ϯ�<~0cב�Y�� �B�90d62k�D��m�\�:����j�@��|C`��J:3[+%��W�~�c�2��Bl �Ksj�#��$�)0���r���:l��HI�pS�k��WHw���4Z�ɘ��p�Q(�n��n��3��-�m���E���S6BG�E��^�F䷸��=���&A��=�=bΞ��E!^�6B	�8�5yѻ|=���y�c���&=V�.���}WL.� ��A����\��߀��,�����2�}/����{����r"�� ߽u��-�_�k@��ػtoR��8V�XZ��l1��.Ԡ�1��\[EJ���~���hB���y4ȳ`j~r�h��
�h��g�߂�|�N����f[r2ܑN��q������K�E �d�PmW�4ʉE�P�L�0�_�%H��<H�ua���M&��C
�G�p>��h�.��`$ߑ�G����J�,�G�_G����N���oS:�@��Q��k���-Z% �c�}� �4��ۗ���#p:&-7�V3Ƨ��]���.��X���1iE~����p�q�G3�7���H\��CF�_�kҼٱ�댌�הtE�-��w����؛���.���z\��S5�{um�fump)�=t6W�ӭ,N�c$���$>���[�/О ^�b����;�������b�
�F�h`[(�c�m��{����ւ�@��AqCx����{G�J1ď��*+�����t�37����O.U�=�C�Mk�Iݖ��!?���+o�~NP.j�p�V�Hk��%��?O�)a��^&ÿEe��1��GV������Z&r��nOZ�7��B��E힝�NS�ᵌMe�cN#���K�)��9S�H=�p�6��#mL��5/���b�@�|��˦�-��5�T����id�ٝK{mK��-6O����;/���"�3BZ�䂄��,Xe��-	�I� v���ù�q�5���HS�0����h۠֓!=�_jĒQ�F#U���b��.����|$<�B	s���n��ݿ�]Ɩ����}j_=�DӮ�~����M5��d����j�����Wt|���q�e3=�����@ô�ظ��	8	"79�`��SD�]�}�O£��&�Ѹ�e`=����v�����i�a���ͷp8�^\+ȍjla0��o#�'�)Q�<��t�����]��r�?��J�{��B�	sJtߊ�(+A�y�y�Fz��,M:�kLXW8����-�!^��Ok���U���픈�T�p��ᑅ�:���Y�%�L���T����hJ��*��e#���\_U����2���7f(d�?Q�ۼ�$��|��۴�c��R���d0��k�� {�Y�Ǉ����/;��W�A8��>~�+Y�����5gP��̞2���D��im˾����F�\8(`U�}�7iï� gt�E.4�7�Os1z��nͯ �X"{
�ɸ���n?#5�c��,�~�p�!{%�5�� X�� ��m�:�I�?@>�eG��J���mΟ��Gx�A?ίba�� �Ĕvf���mO{m�/��[�r��-�Oe��E~B1�? y@�	��'B�G}kw�wM����}�����Y�|��Q��(҉2��ΣwZ����:r�ޘ���K"yev�Qp���#T�0��WϨ�h=�~��2�D�ZK��PT�B�#�X*��"v1$�؍/hh�T�6��A��WM����Y��a�3�OKY�E��̒�~���(�a`��e�X�~���p�����J�2#�z@
2;�+͈0�;˵ �IA��
��X�����2����B D�D�M�b�ss�Q�1/=����Cp?�K���pe��M�����5�|�O�����
:�Ϡ�w]&�s����i�t�SD�P���F:���eck0J����'V��/)ǎDjx7*a�Wµ�L{*�z�'P̉.�M�A�>�Anh��d����a�i-��b�?q:˖8��ɟϘC�_�`�Q9VԾ���yˢ�8�)9MT[�) T+�LEŸ��j0�ɷ���ɿ������a����t[C��	���&��Y��]ջ=����
�ł8!�(N/��Jku-/C�j�)ڊ����x���0��۶!m�Vr+�ʦFoY�n�	��go+9ǅ�R����\	w��J�ͺv�Z����M���hIl��@fs�s�fH�Q�����<����c��je6<��u���5c�8��,�,|,E�3s��{�9���nŊ��ޫ|�����#moc}��r8�=������f�>���v�?${}�n��O�<DvK�h�:'�+��Vr��~�zň�"�&��8M�ƺޞ��7I Tt��<!te����݀吵:�ئ]�m8�/����������Y�j��)喳.�و�N���j+Է&#��|��7���c������v��s���7��!Ӕ�J���bR�,���=,L+��� iu��g�4�h��Htqo&�p��t��0|H~�U�H�1���U�|�v4t���l��S^�)��ʅ�m�<�p�&t�gRQ`v�sG����6�c� A<����N�MG�I��>��[�O������@� �oKJy��-�|&���-�N�SB��,�7	�cG=�g��i����Ð�N����h���xH�eb�s�[8��֤B�=r���b)�v���T���[�n��s�6g��8�6��q#&�o7��� �S'0�?����7��w�G�<u���?sx���3�hؽ�2�*���������j̯z��;�YxG�akr���WȼD����jm�����Fm֫:�d���+�
��\�=�r��d���I�*V�ࣄOE��0�yb4�:�g}b�BQ���z����c3�;��|�e�L�v���X�W���?N�)��!+"I���9f�~�>[��p����G���R�{K!w�hOs�St�w��H*lM����k�Ӑ&z���/�!-����',�wv������ �������vN�&�M�����몪�����z���#��s���]�ԅ��nn�}c[g�y��!&���Q&;$|گE�rC��� ����|]*&��h��5 ���Y9'IӚ	��-�1\�<��bN�Qk*;�~(�̄]U���k	c��^�]=*�Nn���w`�g�\��n�a�R�"����^i����\�9UK��O�{�/H_�"J�;���UP�ݤjXS?q~;��1	�x�x-���ޢN�І���ǡ�'_�V��jg�(^�TrBaT�-.>O�֖`�9�j�h6��Cl�
�_���+����@��HX�ȟ�����1>P9��=����MO��g�#aF��	�eҔ���T���(� �Mk�4�HE�����@&���KG��,�G,p��gI�@ ��	�Q��:?��ͽ}~$sb�Ԏq�!p�5�$a��)�@[)�*����+�q�[���BXR���\?��i��ck�ڴg�%�#�����Fx˞���N֫:�N�����; �+u�ᾳ��7I��6K�wAO<���jm$�J���ۦ���WS�l���>��(��F.꿠�7��b�	^q���pi��k,䪱g��T 'ƛ`�Z�H�F+�7 =VX���@g e�J��}[_��:n��i녵���Mw-������+����Ee	(�v�ȞZ���W�L�,r��T�c���@�����)|g��C ʂ�{��#x�+k�ү��.N�t�N����S����7T�e 򅳲m�'�lae9SҶ�G�k*`�n枉��S���E"�T�����S�Q�!� =(i�4�'��~\��a��@6��?�X�v�^95�a�����r���_X����=�
6L�cx�^̝���f��^��Θ�w�'/
L��ڢܵf��'��!�P���i�]F�>������HԤ�BI��ȕ�"H�P|��T����.�	cB+���l�'W�q�[	5^���r#j�G�;[F}�>����u\��6E�������#���|ш�V`R����=ŒIc�>n�_ [W�i��9U?G@��E^���#����BJ�vL��s���u�̞3�E5�Mf�CؤPa�b#g	<��̲��~1���G����)'}C=�� �z@�3��R/� %�w�qy:�sw� ]��� �9��.I�4�^��U��C����g6ێN�v��<]��W��x�!��t0;�[�G����{�����#Z��##0Sn�0z��ϓ��;�t8�ļ/�&<�fX� |E���K-�^��#0����-y��h��i$��G��KRy66�mG��:�Tk�0�q�o�`v'��lS��u��a�F��l�¼2c��1��������h����I�Lj�4,�. ��,��ϑ�[ G�]Et"WD�)�{��N��}&��2�;y� ���հ,���+ � �\��{Y���O7)��r
���mȵۯk"���ձ��*f[����ئ�-=+���<�!�Ũ�R���}�`C���h�]dli�o�̥�Kw�����ո�������;P���N-0䙳�d�pZ=@ؔ���S\�!�hy����i���R�f�R��]`�@Z�`}&�z*.�k����{�V�;�|Gj�R�z[�3c��M��Y�T8I<L��i��KLܐ����U�F����IA���|WOf�;x����z��T���;��"����$��#y2��n �}�j��!�-K�8��g����.�M5����[�<����Y@e���-L�x^_9~�E�C�WG{_-m��M[HH��1��9dv��x�7Xb�뷙���/_���m�����I��Y�^��tp�,/����6���q��Z�^;"sz�yTԄ���g�2��<�2��x���?����-[�JW̱5g�����E��{��n��D"mʁ�cma~@z�� ��Zb��QBfqs#/���_�f����'63��+�[s�jpe�&R|�YHޏ�N!!�>�I��1�ع����_��0a�3���agg��i�Z���&0V�+>*�6
�k�Nεzf�n��v�sqa����Y�:��3��N�9gN���ua�{X������@���VZ�4�Ɠ6_�r�JIʗ>T�к�A��r'M5�J�@M��d��F��H;�m~��8��iI�l�_9-v��ZҘ���!(�Y�i����]�|ճ3Z�ɉ�� �|������r��W1VV�_6�,d[�&uhG5poo؂�@ru� s��v�d>9jN ��w-r}܌�#���&������_͸��u\��r��A��R��������%�[�F\��5��7�پu���"B3F��7ĒE��<�(�Ikl���N�I\)���Їr���@웷Ћ�z���MX��"ې%��?xfc����Q�bN�b����8l%���=��Kv-�xщ|e�}v��.���=���6m$��.��]2�o<^�~�R��2�IY~�0��Hcm>�,�g���;�1
Q�:�D��N�d��j�����o{���Jc��Q6v^��ld�%"B�3��}j����4~��V��·[N"5�z����_�n��RDʄs��~�aS�']z�-�N�>�w־}\^ �kG����@q6���I��qO�_���s�'���m���Xuqk���+�jY��*Z�4BU}�������$/GBI���i7k����_����G�Z����9�s��8dY����	�.O�>��:�-��F��� m�!���n���m�U)���8�$͊�'�.e�xH�4����f�9`<�M5rr�F����
����3���"�e�,%ؚ(gtg8����H�y0j�o]�U�@=cu��nim�O1��"CO�5�٬Z�N�㚅�L���Y$,�.}A���6�R���B��|�<�k�h:�&��k~s��i�s
�D���[���fvi`#z
&7���n�ݽR��$Wv�-���(h�	k�N)j�p>�d��+���c�^��N%͋;�5rFn�b�P}� �D\7Ż�-t�%���mޓqU@g���Q;�qo.v&3[>�G-o����ƌƟU��ز�pg,I�Q����>?�`��p����Z]��R8a�!��������׏��k#|@}�s�{zMV�u�蛣+(�3��s}�T�'�d�G��N`eT������X��$��z��d�5�$���>X�C>rz*7��)�*y󱄻K2r����ëP�rcJ���@�HR�9�=�;��U������߾Zj���G K+'�z��G���:�S�g��:��������񼼼�#�\���or}�nK���'����-�s۶}��~=�ə���&���h��ɀj�?X��ad"�n�	]m�&dV�o!��Ͼ#l@.1�?���:J����m���
���~M[U���n��/�@IS��tl�m��(I��\b��P(k]�W,u�(�:m��¯ؘ]v �G@��B��ӻ�غ���b�U��(�R짳�l1nEP�$�^��	툸��Z0\nBm���	޴f~���t�c�P�i$����P�xu� 9Ľ�-�j�B��(���ʾq4��O36N�m����-v�F&��"�c���ՌY�5�<��<���e�� t����->h�}WXN�c�o6�l��Ø6���ʒ�����8r:�ՙ��N����~s�
��bϚ�/m8p��ҵ0x<�ޔ����<�]Y��P~�	��o�cN��4����c����Y4+�"�iu��O�DV��n?�����Q��q"��tћ�֞�M�̨Q�~(C��Íl�#���-|��p�cQ!�IyB�5�`���3S��8iU���n���o�_?!-�>"�?�(�~/y.�:D2��<kǘY�	!O��w}{2���X�h��gA��@���,ʙX!�ݱ���4�ȧ��it�����)�8(�Z��f�[��ԃ	�л����\=���P�3�m��ѵ1��J�Ϳ�D��Ұn�=��1��x�}9�#=@&��Th�a��(������A)����%�!X�������X��-7��V�Yȱ�}�4岆��'!���J�ێ��}K³l���SN4fdH��q&mU���IG��hOv_�o�hH8f��^Z~Ҁ!/���һ��n�${�������}H˹�i].�TtB��hW EL�'�>��׆%��s��f(�I�b~�em1m@| �u������K�� �e���v�-�eE�"��U�={6(Q��h��ćw�r���Mr2<G���H�ٔ8�X̭g���"�Ϩ$��BRE=�7]��@� n%Q��&�qJ=E��}�n7S�w��=-U��6o+;9�8�Vא�vϿ���*�|0Tx�d�X�
m����t�E�և @d�w�H�l��=P���Ĝv�����X F]Ct�C}�����I�� |������⊳+pHx��"]n�+�?�k�.K�"�nhk��~��N5��7<Mz�P�Ů�/����Zk+(�j>��O{�:�"�!���e �h9�S�SP2�˶A}x�\�Ͼ�F�����v���I�>�0�Z���8zU�䃢���6���2Y�#��}���ȳ�������s�^��}������z/�5@�4z(��쉤-z�u�#|�>zmȠ�r��o�*j�w��8)��ə�������猣hO`���/Oʫ���N�"�E(b��2B��]#=L��+h$�2	�2r�:wW�xex���H��^��A����2�������z{;��#���$o���T�T� �;��B�Z��/{�z�)�Y��ߚF�3]&p��#���O������{W
�P��(l�h��.��/����V=A�{����[�?��=".��kڽlVM�c����vB���\�Ib�:�� 
����S��r�	�f�7($��[z$�f͕a�u&�r�FѶ���SJRp	=&6�~��D6�s}����>�r~}�(Ǆ�F,�N�k�c���h��k2Ͻ�[�P��g�Z�9	@�i|��O��#�wi����Y��bX�&�w1WI�i(('ن -9��9kإ��[ܯ�W��V�V�Ǫ�>lk��k"Fz�ؒ4\��$��
/?l��$����F+�!�����Y?�{�K5w�Ua: �^�����p۱�C1�?F�w�7��k���c�~��)<���vv/�U罫�o}���'��;]n��ーN����5��6�`7���u�B�(�!:�UO"�������ѪT�<ws ��9/Tg�5�g&��ag�ojU���ά�L{��=�ށ-�8���B:�疌5 ��S쏜���~��%"��*r�L����祿Z@��J�M(�
E��d��Ę�"����ro��Vh��QhҸ��F�lVƓ�o��{.k
�Qy�sx�h��3�Tc厎�߷wl-L{�0?�?�P�qjb��%�&�\'����TG�<aa4���$��U0�|-���� �u��/s[�ҳ�aa�p���8�H�S{�?���{���!#��/ EŻ���R'�9��0��e��ݾ�Y �'W/k�^�_Άe��#$@L�I\R�>�ЄH�u�Y �-�bv�&2�׎
�9�棃D<��vY�{�>��q�Z)G�j��] w�3cCH�킑�vWG+��xJ����j�����y?��W�ԏ83���t���ܩy�?{�YI:58��>�KĤ�'�<ڢJ+h��RJq�߯#g���M�m���^o��߶��Kh��=E��p��d6r	���z����H{m�K��Ӓ��h��y�*R
��&O j_�T��c�H��=zY Y�I��7�T��klL�4�;t�0��G�lbۡzo�ngj��%��w����v�!/�S�P���ZcNT'{��l�tC�l{�s@�n����?�o���na�b˂��(�|�bbJ�+=��'�`@���R�@:Z�{���������I+ ��@������߻ڊ���n(��_�Z�F���%j��m;X�"<9ژ�K�u&;����Qs[�V�8���\fۢ��-P�mv��t�s63[��#�π�4AC��64ʶwt�l m��~J�õ�,X���p[�&�P7�n�ԩ����fN%��>P�b�����r��+��{���Y[*�jm?ۜ��T@�v*	A�����$���7H���uz���$��� ��<'������y�y�42'Ӡ��ʄͶ�~EhĊ������s���F�Jj~���B�C�tAW"�i;��l�ݗ�0�G/�����1|T�V��	�OW��~V��涧'�fA�,�$�0����7H��>�(~N��w�.�-yYO�6��D ��;<���{oO>���0�+�'��ч��l��ZF��hQ���8����(.��n+a���eѫ~�Ak�0�q#|	�0T�
�c�����|��B��x9W�c~*)�r�����Z'G}���o^z!S0���r@���?���'ew+�����$?�q3�qZ�������F��^A�y3�@�����2+����Rb�{�6�J�?�j���t�!���B�dO�X1�7΅�4�M��{���!��Y��5�� �,1�%v�8���T�pf���U�uTQ