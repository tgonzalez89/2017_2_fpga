��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,h���~�G��G�j�V,=�ԸL7���[��"���:mL�^����������?�ع+>�M�.�Ih��X�.�G^0*�շ��د	��H봍YZF�l5&�H�a�q��$��pk�5A��n]wEp�J�d&w�)ތ���k�9��p0�N�z5:�+
Y�(�K��?֩�2�/EO89O�Ѻz}���I����&<��̃��$Hŝ;Q��rB�+�e\����ԺI(��;��5�*4�X�I ���U���c��d��W��X��%������l8Ϝ�K��_\�pM�����Ű�Fk!%��)�B��mV�z�g[��I�c�VY�F�v��>s�#O׸��6)O��E56#6*%�����K���K*�R-!�6`���f��Ļ�C�EA�S��`�ٰ���w��;��(͂\�{רS<�s7�����h�_lhH��r#8�s&@<�,�ݚ~��!w�M��m�P^�ʂ�Z�/pX�1W�,e����x]��7h�������n�H/��A���e;�5���J5��k-�����:H��$LjNv��?j8�ߏ�gp��&3��A�"V�᪷�W�I�E>8��kl7a����� �>���,'��)P�Y6�TX���z�"��"sDa�e8@���m�&ٔ�k�V��˂��gK/D|���� ���{��7�����Ā�UK�&�?9�+����<\aR��+^&[��È^b��,�}X~>H6�s�����V*y�N#�CH'Z�`��x�J����|r$sƜ�=v�s�@��:�������,H�y:B5���/��ͺ��
(�xho����渓2S3o��=��'���������RdqA=����U��h���JR: �TI^�O�;�JuajH�x���<`o_3�p���U���$�yb�K��^h����I��O�,�̛��;F��ix_�Nn"�:�x�p��&�w��̚:�g�U{��=��~����t`i�phe��ԛ�*�
���=M$��%x�u�!CI���)b��u2�2ȧe�%$/�;F���q�3���eQo��Qk�@�xl��j��qs,P W�A`��'W~�����F\��/Ǥ=Ф���[z�U[Qa���;��N��Lo}\�Уީ�)�&���KS��%�U��?��={��֋./s��y�;��ZK$�{�žn��8���x�f`<�sV|�;���GY���MKUg�`z�'VIV�=#L�09��͸���&� �7���i�X��'�c�( �i��#�՟�oI�R���|/r����9`�[�hu�=P�0� ���5 sY�4#Dw+�T�D�{�}�f+ו:�-Y�eⳟ�`Z���nޅu���D8Nܙ��s��p�3��b�tb�V!��iz�i'wz^@L�ϩ��B쬰j�Z��l!eyR�H�_���3��<03�~�%�.�����**	�AtmX I�>��?�Ch���%��ytu <��H�W|\�ݭ������j��B`H���j����s�D]q�R~	����A�mjp����X�妥��84 �zҺ[C�QRK�P��$@�&q��OĠ�O�����\ӦZ��JY
,�g�\0fŬL����sI��Y̺�陼!���x6E�xZ�*4N�#��]ּ!�k�P�"�%j�ᝅ�P��%T�E̗�,vW����ڔ�y�o���.�Aa�"�w�pC��Dwu+����\-���W�p�C+�P�>Y��}�������&�Kné�i�|Q[J�� C(P�h�I�eNPά�s��s�k���*����&�$�\������P��iţC�w]#���v��b���%�f���k���+=�׌n�D�T$�n��&P]=PNz�O�u����s@�}Z��vr-��Kq0g����Nr2���X�Q���5��#�|��K���m���U�-��_�߰���*!�ˊɹ���1��{Úڸ񙹵g����`��{���3�ESS�ò�HwE���?�0F؆a���Pn�i�6���CB����L+ �gq�=���:J3���-g������7�jU[r�����*/j��0�$���~a�{��Q�%X�d%EZ�����S2�ғ�9�l����C���$^lK�W�Ԗ��FZK��?�e ��7L��gO�����/�5�T�_^x��.�(���0�7ڲƏ��Ѝ5��&��S������}�_Y�B[b����QcWT%�4�����هo�C�r���?^}�cg���I���|�[cȵ�I�B���K��z���jr�{�%�C��g�ѣ���'k�"o��U�+,��������՚wN����!)w��L����gZQ��&��syi��{�Q8�>z�J�u)u�U\�'�v��Zek�.�HO.��H|4�
�9=�p�h���e��F M@m"(˒�0b;�/��z�F�=��d0TJ�'N

n���??P��,?!��H�e��]�Z@�ٿBڠ�!����Z{[��ϻ�`���}"�9�+G'��ۊ��A�%��{�f�I���Td�-кQxr�`�	���Q$���T��XxOl��>x|���#�u�*Ľ����r�������+�B6'�K�K��X����#*��D�O<�ڸB�&��2�����tG��8�AN�:�'�+8��0&�7����"BV߫�y��]�<p�|%�ޭ����u�z"p^�I~ט����5�>/8�N��SW���+�Ĺ�t�J0����.g_��CЃ$x`4:����pVK�{�>�r�9�>ox�ϣ�dO�{4eiq�l��rɎ�qT�iꅐ�� �k�7�Y勫�BoЉ�;�w��J��u����"pRnT�5�n�m���m�p�I�}$�f������\������V5A|?�Y���é��z�q����G��3H�+����8r�b�BUE���CE�mQ�Z��x�
_�yg���%�V�M�y.n��9�c�H}���Q�|Ǘ~�����]&Y.	�h�H:Bl�*��bn���	g
�O��ݣ�kF�z#0g�,u�&�n�n��X�	�ڇ����=�*;xP�9������z�B���l; �t߁�}E��]��M�.��0ÐR��p�8��c���B�G{;柯��ϚW<��A�Nf I|�&�,Q-{�K�R4��L����u�@��w��^
 �R
��n���?����q���f����������kY�yB2w�{N���*E�ݩI]�"��c:�m���&�e��b�M7A�Ӑ,gҜ&��e�Uň(t�k���q�؏�
��|?D����}5��ū	�����%*��s�'�����������{�
y�+V�A���B�_��b��۔�T��l�,���$��?�E��Qd>C�m�q����̧�������?+u ë����1��)VV�2�c�HŔ�G`\(��/��0]C�F0h�u,�7B00���~�`.��K:�|[(�.#o�$� T
��wv�*'�^��PȤв�z#ETMf{K��BD��;���w��.�U�l��Š�D�y�k+�{�MO�
�_c!�/j���B#p�A�/�<zw�l�}���l4KSI�Q=?M4B�(�p�\7U~9T���}�S�a΀�6�8�y�Ռ�]�I=����V�1"$ѷ����yP`g��J��M��ˆ�M}����_j���3��f�s��p������<7xbHI�P=�'�����2��?�'weE������j��0E�x������>&"h��+��Zn�O<.Jt�@@��?�3�@ /�K�SBQ�T$K�������߽��*�?����r��Km��Vz���z�A�o�-&����-`�C}�_�y�Z��8�.��W�L����R�*)�g[_���T�}���H9��%/ū�~�21+�")R�F�%��w-���:����vJ�_��_;o��!���dŏ�I}dfv�m��0�$Ʌ��7&��������5���7�:��s�����*��+�DwkF%��EOَ�jb��~6���f����t֎�FYp�Δ�y�xY5��U�����^ i���?q����96����hb�ZX2�:C-ncT=2�*W�ƕ� ����"�}��cz�����7h�/��±j9�^ǌ�R-q)V��F�BFvi��$��/i8(�q�`a��ɦ��E�_� Z������]�ٴw
���
49p�6)Q��ᅶ�L���lLi苋8H���T�o� ��������:\z�%��+�j����اt/Fy��2w��2�N$��U�Ǿ�Ԧ�`��^�dٓ���I&|�ۏ:x�	ۑ�.��/��N̘ɩBC�G�)Q9��`��K3�1+<s�"�{9�;������1z�m����/�l�GW/j-�4��hWy�Ѵc��Ɋ���&�r�HXr�Ξ鹿m�Xr]�n�4?�e���4_�-���R
�F�WRwǷp�fRs�-F����Ί��[�k�vB�I3�f�Z2�R%A����*�up,�ϭyD�x0X��nR��g�P'���#Y>�3-}�s���szJ�����QM�Y^)/�\��F�y�y̜b�`�����v���<���%���Mi�}�_ܠy�zXn�G�+"d1����mՀ�i����<� ?(��c(��=��]Dk]�'���<HO���{y��<��F��}��b��U�V�;G�=}�C�u���c�Gc�O��o��Vd1��$K�+ˡ��E��ЭM�&;�J��D��ƚc�;�q�N�����:�OL0�|زaq�oEh������g�[�J5�/%h��)*�������'ߍx|;8u��u����ZY^Ɂ�!]q(�85����?F��K�'��6���B� !a��\��6�<��v�����]��Z��3[G�k�����'>�>�Z|���Y7��a���i�2��-> v����I�7ٚg����l�t�bc[C��� �&�l�����}���a��:�ዕ�ԫ��:6yH�x�e1Z�� 61s�A��� ̌:�	`R!�2'���v�{Rnw�9�Ώ����͆U�cB��w+;��f-u��B ���&|u��*c?9�ܮ7���&��xr���@�����w�y�/����=��ӷ+�~��8�>�e����v�v�~E���}��Z���_Z��Kӂ �M��R�[e����G�!���ǁY��N/3m٧�^��6r�D�K�IS�3Y�7OËd_���8�W�s{6��3��\~��R��/Z9(����qS��)�f�����k�&g��Gy47���m����H���-�3�#�"?s/<+~��D�wXg�:ܣ��d��P�SZf��O���� �ͪ�p_�#�]�^�ǔ���t`*l@�P;�2p3��rbS��E"��Pn�V�Ҧ%)}�ߛ��Ȥ'�)L�������R}�X��
�릠:�a��rGp�k��j���	h� �b�V�AC[��}�RT��R�|]�l��p�.U�ֺ���e����!hR�@#I/�R߽�&G�ʫ[-j֦
��<n 2�,������GNC�I'���N?���	�5�j��8�ٵsb�y�ƥ�xj�qm ��	�\-A��a��'��_��ӧ�Z���_%*�Xxٶ)��c�o��%�u��$���\u��,1*®�/fjmS]#Z�4�ܶ����L���RC�_��vu�V�?q�#��q�si.b��Ӥc�� �Zt�Z�ژ��K/�<oc�L$��=��3�N�s�6��b��>���g=�L��`1��	�E�n� �y��+I��53��V�4���%��/u%�7塾j}�{6g~k�Q��p[�Ń�\�[m(;c~�E��~#a��X���3��' �6���HfQ�r�ACo������ ��4{ <����tH��<�!�W���@�����v"�KE�u5JÑd�C�6���ͽaZ���W��7��_����s��T;���l��ț+�;�C���X3�y�z$��Q�@�H{��z�T�e�C��qN�,3~�u*����yJ1G�M����}<�
bK�D�X� �m�Wܥ�}$-���Hvξ:�b�D�~<��h���0HG�"�#�w�-ZA���_0���n�td�2Z�{<a-b�$��y�[>�tBP/X��*V3��xD��ПYS�*>s�#���F�C��əB�V`�J�n����$_�fE�q��a6̅$���L�.�/��ƙS��$��ؙS��qd��V�ʝ~�5��Itb���3f�,��
�h��C���JDW]-��NO�:q��N����C�-:w��/�=ɾ�R8�Β�t��=$Op<�=�W�e�n��.���T`�a223�ɇ�YgVglyd��ԨL����i�������*�hT��U	e�)�&yN��Yj��P�#�Fwv��6T�-��.I|�0��6�2���f�O��]U9�t)�g~��iä16���o�T��گ��iC����)2�Ю4z�e��������x��Hq���|�@m`t�Z5�(���<[њ�1b��|}�e�����Jw�]P�W
D����|����Yf;�=�:���3��S.�ɛJ�- �k�<�e�n�yeI��
��n�0�Z��O�4.�ԫ
�Ea؀��}���܈V�I��8t��]���K�R� �x�)C.~�W��x�-F*��%c���?�BPD�j� ���k(��J�D���î���r���K9��K���YE���ʑ�-�t��-<#��И5�^E����շwTKv�M� >�(}Yv����=����w*��k�D�@ ��������Za�s�R�\��{���T-��)h}a*q+�CB*�U]a�c*7`�zY�
ߌ�K�͚��?k�J���ffw�,Lb6� �qOæwfACA�WgJ��@�P�#Y��&�{$���(hwwb��Mˋ�;>?|�Z�����Ĳ��K���%��iUD@K���=���d~&;�!�F�=��i�)�N)�u���cM@��������ۻ�PEV��x5K�~�b�j��vU�pO�3�ߙ*i��R�x3`�I<T�꧖����#}ڹn��w������
�A�1���SR��&k��xr�(�啹��������21�����'ڜ%��T�0c{A����K�
Ԯ�/~��<�]���	5OO��GF���L�cͦ Kz;=��/��t���\�K!��ڎ4_����~�n��A���Y�E$��lY����`��7���J�ZC,�i�.%��݋��!WGQ>D��,1;El>�¡k��+N�¦Cyq�#�"���cЏ3���&޵�r5�4p��Y��ا�`u+�ѱ3eLV-���泅�*\�gy�mY5
��Pn�ПE��qT�QN��� &o�x�,��^2��P2(��5�'(��{����7����ᭅ.�������rl����pR�G��E#`)���7�%jT_�����4�!���x�2�NZ?FǑ�4�� {��uu��Ȅ�ə$����9�Ǣ1��Mш׾0�/���4���>���霈��~���m]�gu��>��� f"qP��4\ǝ������8�Y���#)��Lyqɐ�dl��b�u��3�������KF�}��Rv�F��<LJ���`�F�@��e���U~?�T��}���9���b�ި��G4֮QG�dN#Kw�z#'���u8S���8�ߩPl��n��0ǻ/H��L�\Q���M�K�#B������(|OP���1�X?)���N5�gK�>!u�6|�8����v/�G �X,a�Ѫ@zV���@�s4�MϹ�4��a�k>m��
���WG1��P�A���i�e��c'�[�"����o^k�<�-��K���D��zQQ.�n��زfq���l)�E��l�#+�����ַ.x kQ�9x�{}:F�	Q����B9��ˈ������*0y���`ojS<,��IGN�%D�:uD!>�w'N"lӈ4�<7�Q��nwԝ��9S�������ͨޚ�}��"�{���J����'��l�=�j!�r�O�S��%=���N�	�j;GHwr�Q٩k����_��UHq>�%R:w���XS�Mʊ�������>��KS]�
:����_��p� a��SgKG�{���][ƃ-i���C�z�� (j7g0�Q@�t F����j���!E��{�o��L��#[ |��.�P���������a��3��y��IPwzT�;��t�BvA�V�J���$�K2�T��ǹ��#-�Z�+!NuG�;n���AF��F�d��f|B��ׂo�`�z�7��|�lT�|�2s`6j���c���F/�����&�g����3N	����'~�-�)���D�]pj"�؋5VH�|*<3V���K!N1�$_f��7��H�ƹn�X��`����
y��A4����,4�f�N�:�M"0W*8������%�Z�P>�����Wn�qt���%��ˏ����3Me��j_IwGr�f6���������%�
t�&���������m"���Y6�E�crt?�����U�'�^�{&��Ӓ�c��,��l\V��3GV�27�@�DPf\�6j1��k�fAdݗO�8��C��9�==���_5����l�v����s=װT#%yl��#�y|�b��kz16�;�S<N"֣�#ZrhŕYE욍�{�y)w�>�i�>�:@[���s����bf�qjpηo]�c�1�
ߐ_�gV|���F�+n�[[��M����24�W��ّQ��.�$[r����kO3�ƍ�;X=�̀aQ��B	��(n��y��ā�y̬�)�/�{k(��3kL���nR��#B�n?�:���f�;v�����,���s�U�����g��h���Ф�V���r�9��u�Y�

��ENVSo+x����3��wd"bH��/&�]3�������]3d���_d݅�:�}�re}�\%N�е����hH����5��~��1�V��c��Ƣ&�����b�ܸK�K��caC��/�ݥ>���]��Z��+��|#�V�}�2]��]ё�P��zW�0͝^Y�MM��w� #sօ��7[�يQh��Twj�׾m��<����e#�i<�FB���းϐ=�]���$���|���=�oQ�t}
$�XY�|N-I�b�L������}��%����Oæ�Ve��p��V����R���x��_�"ǣ�"ݪ1�cMc�}X�#�a;�4��1$���7�~�z'�1�]�(�ak �;reW���N��Q��ܑ؆J�VW f��A�a�.�䫶���a�r<:�%�St�7��[�uHO:����Ȓ.��{��9L��	���e�tN#O�G$��um~�&k�>Bk�`,�n�;�?����|˘+�֙��s77Rig� �~Ѳ(G�5��0�K�������!%�C�2�nD�F>-fG���w�C�mm��hT@����1��P�DGФ�pD(�~���H��PJ���<%�$dۙ�UR�Z��[�
�k���1Q,�LC������5G�i����Q�Q�og��R�9�H�x�}ۥn��r�3R��B2�^OR�C��\S��G ��'d�K�DU����t��E��,4���}�ֽ86t���f�$�Fv��}2��_�^$�h$6>?%�>�Q�l��/�S����\�A��	�jn����4k�i��o�|����Y�p�n���!BׯQ�`U��ʄGͨ�D��8Z�OϷ�Vr0ܦ��9��F��E0�pa3��S�KV%0&���W��Tɞ؀r�nC��d	�;���X�C�v�)h꾸*p�2("B���r��N��{d��
�՚m��V�42�Cs}��x���U�I��M�L��6����E���ly��/K�r>u�[o���lA(��Q�גv��Sa��@c�)�3Ѳ�:9`�"ȷ�k�b��=�|*�� ��K�aM�+��5�Z"�B�� ��3�_-n��.�`�P5�o�Y��r,MU=�;�����j8_�T3{.^��(q+w�[���x�����?Z=� >V��c_ӭX�m۲�&��<|�����׭;�=U+�g�t0�fM�ܔ����p=�9�_�9gb����_��	p�vT�Jjdgpi^w��x����gST^�D�T���E�Ƚ����й�[�M���!���,�O����_w�W'[1vz7KD�F�<5dD]E%�!��!)>�8����|��*��ħ��p�͆��� �>�*�睃�#��"�г6x��5���$�F�=��N�1̥sWǜ�5�O����Zkeu���3ʫN���U��
�Y(�k����oU�w]2�q����QojD��n����^�/���x�o��2�	�QÃhe`���2+��
�BX@�X>��iҺ��5xz���"�a����Nd�~�6 A�˷�y/�f(��KuU݈��b�5��s�I�Se�2�}G���j�W)�2H���y�6����X��t�/�[S2��}��sE_s��.,ւ ��B�n����q5j�w��G�����ߔ�ď�)��ib4H�|t�N�;�ZR��%X.�"uk]�ש��`K�Sre�T l�`U�ϲ�Is�:4�;ނ~�D8߭u�%\
(#�9�q�8ߛ*#���?�+d=pc���;�)��H��(c���D�#���O�_5�Y�F�h�����Gjo�m���p��|4D{���z罁`�+^�׸q���(_m%M=�:��(��?:n
�q�a���	��e�ؕY�d/^g7-��<��xS��S����q���00�E��q�Ո"��x�b��Y2���V]�p�J�?����cx��5|�	|��@Iә�̸-wN9�N-����㥑�:��	�`�ҥ)��zA�?-�C��t�]�h�PL���(��⼎������ �y���U��M-��j'�墟��A?O��4�ԗ�b��J�:Lt�U��+��iR�C�� ��:���"SD9�hp���ߣ��#�XJ��(3W3o�Q�$T(�dQ��n1A$�]�LYA�#�0��c����MGG����ĵ� ǒ����y��k^�����4C�g&^���	��m�A�ٌ�0k�I��/��`�S8�n���\��t ����6�+��)��Z���7%-�d���n{��WR�%�(�����q�����{�y�E���������+�����8W�F]�|�wq��E�R�mV�r3��{ ��!YEz�&���>6
J�e�A���g�V��<N�	n���������d�~�WD�a.��@��� x(? ��f�t�=��ǽ���a�&�����5ȼNՐ�AUM���-8���Ť��4�cA�Z�� �@DӘ�{\Tb���*Y�� pF}W��r����y��[MK�p$�ҽ|V�YX$Έ�n�Mq��e�鼩`��:�a�gf#��RF�O�)��])��4�{���Qsu7��^�T<����j!���B��5g��op�6�-a�M7l
�fkF�D!����R��q��C���@��!.���j/o(�A��\]���rK��:_�.Ⱥ��8������t?!�������NfB�~�4ZR�?�'μw�t-X�m�%�տ���k��Sl6�g���"�"�M�Lg�ڌ��Rq�j,��LG�J�l�� W�<3�F�_�Ȏ/Ql�+�g;� �*���M{���4ײ}�E�O¡>�#��[9S����LKF7�L}  �"ʓf�_!ݯ"!-����l�i`3u��$�p��,o<z����|85�� ��	�H��"�#��H�n	@&h��F.Pm�}�A$}v���VҮ��9����6�7&r�0U�	�A����1���d�oKD:.��W'�R5�"���|�V�2�*�ɝ䧢�ɜNm����P$��Em����-��{t��Ҙ�+�5���js����LR"s_I���ߜ��N�c��љ��Ky���|~�������M"l�T�'���E�-N�f����:*NT�Hn'g������2a/0��Y�3	���wK�z�7\2���Šk%+����ٺ���c\�_BNҊ���;5oq��(	e��p��O _tٺ�{
������|��좢S+J�?K�.Zg<�ꍭ�K�����.;`�2�39?�@�$����a[TSɩ6y+�1eOx��L/}D�fo��T��֑����~^�>�yRI�[#z�#�/�/�mU��거���?'���A������UH��=h<䅩��>c�)}�K�9��Q�u+ڪ0B��pj�p3�H��㊌}�|����|�!��B�#C��S��0���ب��k���"I����}�����R�����C0��/�e�/!�PV�����"|���0eӠ�,�]�n�@T0�m��|��T�ւ��3o>ުAu���E�{oY�L߫���%��_�$UD��~.�N�"���\������V�/�XXwD���YHY����\��g��34;����!��Μ���h̸�|�d�i\
�S��L���_ '�d�p������4�M�*z��o��pdQ�)�,�l��%퉰w�&\�JB��iՂ�Qpԅ#N�;��K�x��zoqn�ÃY0�}~#��8�Dt&$��۪����@m�t�����f��e�����b�,<(� 0�Z0��+y�}� �����V�Y�;�2}���S4ƣ*���_ͯݰ94�]i��X���W��SKLr#�1Љ�˹_�0p`�f�}�u��%5�RR�Cb�����>�,���J�F����Ԫ&V��mIh~����m:��EvPHN�uLg.���
�@Ɛdd*���o��Н'�)Uu�0wjK���~��C�grID�s}=I�4d �q7�g5z=H�LB�X����<ђe<�4�"@�'&~H�ڨ���B�vR&:����'���Ң4b�Z	9���	���Z	dH�Ex����G�U�
B~��>�FB������n��0lg�{�h�M&��d��p<x�������>��ޔΡn~[�V�y�M��O���a7��@�V�l���F���ʒ�Am��yv5Sx�xu���b6��N "ʸ��B Q���"�l���C�l�?�"�v)B5�����3�W�~'�_͙]����T�<�3���ɑ>Os3P�BFq}py��f�C`(x�^o)���o��^���2T��-�-9�8�Z���j�]W�z3i�U~�V��u�zh��ܢ����@�RZ�U:Ù#^IF<�V�v�lf�����Y�Ns��l�|=�Q��Q�+J*�� �6��B�2l��F�U��BG�|P&��͆q���i�	 }�$�%�����V[)Ҙa��J~;�;�"���&��N4�`����a�j��i�E5v����4���`k>5R#��+NP-+�A �]A`:��KeE�xj�Ea�C����!'�"c�9��t�����ZQ��*C*fzqrL���[�f�'��"�6|�F���G���D�U�}M�_�䅑��z�r1��OͦL�#z��lJ�9��<�/��X�m� ����\C~�1W)��A���ׅO�En���( 
 ��
f�<}f�%�E�EW�7���-e4�1Gp�Aa��� A��F1|�~��-U�W��,�n�t�]��,}&���|C�"��'���)�p�Q���2�W��+�0�sFG����Q��X7�hSx��j�bT)7�r��p����L/��G����޸� ��3l��p����3�}�GoB5��j�-�6��b|+�&��n
=���z�04������nF���s����Ɋi�jQn�A�.D��RF�E�4�tU�[�Q�����=p!<��(��h�_KJI���um�Jjr�Ɩ��IS�����J���[ ʙ��I_.o�������˚�1�~ˀJ�;aE�����ƁU���+�,d~��;��t�N�zc��ah����֛���.^��@����Z#1w1��#)��IK�&���YCu��U��K\(�OR��I��:��W��t��wN%��d�w�h�N�� �ؗ�-.�������X�,-�k��6"�� f�m%n�f���S�*��&,vI��k���6�@a�@�;9>F���f�ڢ(�d�Y�F#�E�y�82�t�?��)�CRy�+~���"0�Ӹ�*K-p��>����@�%̸�iV���2}�.l~n9�X��Cm���p�e:�{��	F��ҲX��v�~o����_(�p$�u���s�l���ó"��*�Ϙ��^�,"��1+���kO�ۗd@�����������+I����j�C˂�,�= ��kq��YC���
�����Ik ��!�Cy���a�C<h�����@���f�Z��i'�I-�[m���wdC?վ�u�"F7Wrj����EZ�k�����6y�����v���:Z�o�I7�����71�ek��t�5����ڜ_8�Ҹ`��J8��`QqQ��
�C�\˃��7��~��pnrJ�/�����xέQmkqH�<%���h&�ė��c�J9��� X"DZ�ðl]�KB�4�[�9�8��Ei�̆j�����	)����@X�O����B��y��)	�^�q����P	�gեWp�tm���h#�9��#PX��A����:Z�jC
�����v~�+_�|���`6�O�(,�}0򇰊������Q��}���;��H����t�L��
��x��l])e�O�'��t\&5�Uz�K����A�#l@��N�UG�x�i�o�h�zH���ڱij8���A���ET�&�]�L�o�"��1Z3h��7.9
��D&Kn�=e�$tU�P���*��	�����j����V�Ø�9���΁[�����e58�M�j*�s���K}0�LvUX�ZzZ=%^����[�vM�?��Wv�U������[J"U�P��{�p��.��ݪ��P��>j&|(�Js��I�op1D���L7���s3/�O.�pDYF#�!�O&�O�@��܇$% ��q�a��b��hNce�p��?Fuѧ
�����D(�M��;�G�p��A��X���à��8ÅA/��Z���bF1]�l�%�x�,�h ��"=�zJ�G��I��٥Wwbg���<���y,����L)��j���pu���:�C1$�0��Z�㙕�m;��C�������S�W�Z��_��[E4���p�
mD$�%�.8��qr�<4v����IW]���j�<���y���>�v�WZ�|u�1����_}���>vp�w'�=>�T�4��h}�SFEwѤ�L��0A�}�Ҏ%؀��e`�ү��5p�4v�����1�)"��`��氅$I�In&��ms1����P����-�"h�y�r�n�D�����ݒ��E]~��H%�(�#�Q֞4��µq�D����O�+`�Q� ��NH�N09�΍��W�;?��@�����Ø V�C`h"/v���8v/��k&)U�1��o5��޼�Y1��4�~rĸP�fOtnu5{���U���|ᓘ�!Aÿylχ�g��tT��?��~�������8	�E�kb��	� �L��7�ĕ�1�8~Ȕi�ZE�M} ү�Z>�0��B�.^�<B�L;�>���.Ԅ[܂���W�:�J/�T�$�.�7o��Z��#'7Fu}�#fï|J��{µ3� gvh����~��1>��M�ćmL Ԫ|�7ӊ���-&�04_A1����[�%&wo��w�g2�m�pGM�"oJ�{ukE�c��ŉ��e'i���I6tKL�e�'���eC�r���Xk��HMw����G����u��MiJ��k�G0b��GF�x��[�u������F�Qf]6^�#����W�c�Kd�=&��}8u=��SƂZuT��d�?m�� �dh����3���� �s�@@֪%���x���r�����|���qPč�I|�7-�U��j�/Q�����ɳ�k����q�v
EH��$p�e���|�<�<�/~�)&��Lr �"C��}uH@fq���R.�Нݯd�euhg��?Jfw	G���������_S����=p?}/q��D�HEc��B�.du�3��$ӢӒ�5+�T��)g�D��[y�¶8��}�����d]�ϩ�kl޸��������J��b�3��_ &���݁U���;���e5Vq%�Г+e`ņ��۝f�|اC|�Y®s��r�+n�T�vzÙ��g������ύ]y7\�j���Q�:y�����8@#�F�*�}Ad�D���F���N��Y?�n�ז�u�^̦:�%��O�@ς���D�T�8+���08>����:��#�}��Ǿ�&�I��=A昌�e���L��v��t���q�X>��̍f4�P�*�{k�fU�-��N\����F�9 (�,N�V��H�Zrqeą6�{n�d���c	ꆫڌNI_-�� �`x0�F���$�%��TR9�/�D�~��w>U4j�sh�a�
�lV��C�\��=9�A�A�{���[�L�#k�*���t�0SG��d�]��L	��hO�jFk��1F&k�Y�7u��F��7(B�"�.?�s�E�j��5�W`���J��;��t����DLCsgȶ�ZקP-w�u�k��UP��u ��eМC�g��,��T����9'�Rq���d�1!����;��������F �V!$xI���E��m���V�����P�Vș��a�� .~�\�9BGͫtg�쁵A�.kX��0���i,"U�n&';JC����8y���L��֩\<�g���4��X\�q�
�PN^�4��I���r���'=ҁ�q;`|^��Ype��m}L+
�0�Y�SL���̕�i�X��Ly1kF���"��4��ms��f�w�XT��� �lw��b�"6��C[)�H�cj��c�q���b��뷬a�07'�٨�Bw�kk_�N6O�$����V�� ~�$[ߙH(aH]�ON@ƏnI]�����K�%Y[��F霏H�3:e�.bj���2ߴ�L�єrj>�8a;�Y.������(���W�ڙ,he��\��e="��O�-d].|���f�K}_{���.��Y}4�ż�΅˧Wݫ��ǜ!�� ��M����Ka�Vt�d:�縃d��cWR�g��z�R�����B��u��K��\�N�~�1�h�xq��U�D����R��%��򌷶~�L<��n�*jya��(�ˣ#���$�"2��i
��{��D:+�E�`vP�?I"��'!�j�����[�LЪ y�f�u�p!���4A����5,=�C<;L��`q\y(��O�GD�y����HfQ�¡}�;����'�[���>�������3Cf]}��p�������I-�s/�'l����,�6%ͧ��a�%�k����6jq��EW9W��9U��0�!�Z�� ��N�����[+����7$6"���8�B����?��|x��7�۪�|�CY@������n�'�
!�V���p�-�Azp� ��Y}$H�zA魷�ݼ(uJe7��l�ڀ�}v�5w��oY���2{	.�.I�.|�J�uW�0�`G���Ѱ Ʌ�K��4��!�|�ը�!�,W3�}�@b�����<M�[Y�(|c�Q�{ٵo|�H��5��f �D�%�֬U��S�����P�< 8�	��laB_������{��qx�����}�k��h�J��	�靵��'��L�Y,p�mDY:cO�Y�ӟ?b�G0�Z��z���9��С-���6P��v$*C�hԿ���"�̟���t��v��1w��:�h*zVЏ�i�噄]ׂ��]�P
Ԁ2�i�J�k��k�a���P���f	�i����+r�06s3���0t�)��`��z�ORʼ���n�jK4���y�B f���'2~ �{H�bj(Ԩxi�T�*@����Hɷ�*R�q�r5��z��a�w��
���tD��vHfZs��d{ֈ��*a%^��j�O�z���ø`��2Yrv¾�H	e������ޑ��gQ(ɓ�.'j�P�.Rik��ݚ������~��ڻ��֖�F}n��Q�����w�	���ȾHEe�{�1���ۈG$�w#�c�j����z|~|s�I���^�,�Y�%+O�u�+>~`o<�Se�~�T� ^At&kk%�����d��~|��2vNt���T8!&I�xY؛Uk=�\i|u�d����.��k��[�9>����(>o'1�[o�J�������6��Y���/�<ʛ^��2���*�?M7��_gme޲<i��ScL�K�Z\��P���i�?�ns��dov�Tӹ=Ю�=��@,c�\Uq}w�kM�ڱ-���J����T���뫥-��pS�b��=�}�7�8�!�5R�[K�f �𸨅�;�Ǌ��ˁ��2��Q�,�I־�RT�`�:��Y����&F���ABL�(ZP;H)�}x���eK�8 D}�5jؼ�t�e��-Z�uyNn�O�|���ЯU�A0�4݇�iD>�v(z{�g��jv��:$���l4Gv'g���Z���߫m3E6v0���O��t����T%گ^&��{��j���}�A���H
�t�����5�NhR	���q�+u��Q�TT��L�_b^��yO���Z2�q"-��l�r�{�}~Ԟ$�Y�2;������Re��2���5��hL~���}"�d%6rvΖH��H^�6V�e`n��ΐ������̥�X�6�	�b5�!���'f�	 "|L!���J��UW�������� l���R6T���=iPc�OS�� �iKI�/�$S�T�����˅�œ�o)սB���5��i��D�����"*y�����ثXP"�J��%.;��s~�"���9�%�IżA���U�����!n�z��A��E�)�=\T"��m��~��TkN$ae<�,.����#?��fi��lI���Ĺ�}�_@"�q�sUXHx�1�}������H�n���ꐰ*�dM��嬕(���3�%I_�rp�]6@�UsF���Wӂ&����Œ��CJ�	S�� ;t�	X�>��o����Ӊ20�ۘ��hA��7f�/Ʉ�2�R`�0��|�<�ڐ���������m���9j�p��T��4�c�	e����,5��4M�'+��\�pE\D4�[>��t�2c�3���m��COm�b�:q��GU�M�e�:�q���H�G�V	�ƹ{��!��� ���DV��C��B�xO�B��Q��ŉL�yb�]�i�ϵ�0�>r>F��n�̦�ڱ�� FA<�����䣤3S��-4P�=9K8�����8�آd��Wr���t�����O%;�D�_������D2�!�t5�A�6]R�L7��.�0��mf�4���%i�ާ�jb�O�6�	�CБ>�`�j͆��>�A�la�s�R�KiQE(+�!Y���r�"	�&�/��:ʙV���V���|ܬ���+SIMl�␀Z�!fTi��4n7ㇷ���ߕ*�<:��s�`��0��?��y>6	e����z�
��OI�Ɨ|�B5aٿ���Sա3[R���ʂ:U�2��A4�A��1�� ��rzUu�Jx0����2����/���t���z97�<�ᓬ�`|�P�>�;��u���2L�D� �+�-��ru/��E�O��$��5�0�$$�2�'�#�y�p�t�!��,�<}���Y����q��2�0|��j�aٻ�a	
���>-A�x��3�cv��Ho_2����z��t�@N�ܦ��囯SD֍Z�WM�'Bi��A�n�@�/	\��&�cT+�9�*(Y�a��JÎ<��R�
\n���6˔�>���x��mE�d���ZyMw;O�rL�?������f�B�,3�Cl�:��5
7���Vzv�4O~�UL}ݎ�\|�����8�nC�BdlJ���T�����K���a�z-8��X"���I،�%�
���D��O�.B�|[#�id�ͫ���p$����4��|��$�!+
C���Ϣ���5�S8B������#��%a��ԓ'a	^��eE�0��L��ɒ.A��a��kT0-����l�?�k{u��G]?Dkb&�S���2�ct'_~���xC��\��&���m�9>!g��1�Gpk�/�o.A͏Ȣ�1�&�5#Ѳ���x�}ױ�H��G�2��yu�D�c�n뫧�Q����Dm���o������"�4E���~ώ�i~T�+�X(���t`�,�==-�[�,>1��O������'��J�rrUK[嚭Sr�4��㲔�뇄�v�.�o�%3���O��cM�|Ww�f �������Z �;�T��c�U�I���:��^�M�r$�ǫK����d#���d�#V����4� z�=1[݂��7�EIK�� H����.^�dz���>s��f�s���u��%�ei���զ��@�A�\Ӌ:9�qQɇW����)y $���H��6!���~Q�4p{�3���A����7}���<~�����,�?���̼U���h�L<��@(#�D@	~��aOVHț�zb�ؑ��b{��'��\�OǸ���EN�hp��Ǯ��*]Z?���\M���N+n�q3�Y��%gb� ���k�xs�&�ZkJ�͜���(��|�=&Ml`9F�Ǚs/����T�s�|����L���0	�끎���|v�k�s�7tnL��6�u�Ը���`!0[��9�:*
�:��w'��ӛT��-��G_\�
����@�)_���@T*�4[����V�VQK73�H�O���BA���D�?ٯ��.[E�IJ��%��AF�����Q��aJ�7Ojz����m
�x^���iq��!tꆇ�~�K��o&������/��Z��ss-�*��Q��Ӂ�&�������b�ƵЋX9��n�Y�!�T
c�W�W=�L�G����CvU>U�Z�'�m> k!��JܒU#+�0�O������~&����i�G�+��&�9=8�г�V΄V��U�IM�6�9�4e%�-�A�o���s|Ș�O��ҍ�}�A���VOڱ�}�0�#���A��̪\Hb��#}O2��o!s;��UJ��.7��p;Y�Je�5���ͶV�}g?�a�G����W*���e��3���J�����{�&�ՐTe��Ƕ\�fo+2W�5�w�s��n�ގ�D#cE����u�>j|�l̬V�ʗ:`�Sy�V�Y���e��	C�Q>�u�Yv���)�b3��˪-l�Ng�6�5R���ě-fgFO�b:��AL�7�@O9�����B��:rӳ�2�N�m�ͬ嗋�����0��6ׂ#�רTO-���A|��T~���?��J��6"g�2`̄Z����g�� $�;O��~�!��i9���>�s*rMwl]B��_�g��@�t>��s��:�P�C?sm���!u���ϲ1�Nt��TtP�O�H-A����>����hQZ�8���<�j�s��CIᜂ!Q��oq�ڿ�2 sC�FJ������.��p��9+LW��7�`��x�E+
�3����0�&C3�����UE&B�!�(A��U�&;��TX�ysx3����^�<�m[��Y���ˏ�Q��
ڗ
mC8�"9�}��~+�GO�
�0���i�e9؝x7�,�M(���OV7�^�9$�M���G���u�����5�d���#�☂�T��Y��ҩ�>ҋ��ݍ���7K�MQ�ҟM�W�l��H��%G����&]ޝ��.ar���h�6�Ս�D:A�c�r�G.�#�Z��y��=TKT�Nð�B}��s[>ZgK�,������+��Ow�k��(X�٘y$��m �!	q�}�,�R'h�]�+�7Ib�ӴDy�D���3~?��� u�!�Aa�*cC�/�V���'@�Lȕ�^V�P���'Z�������\z�,�	�6��h����"=L�!�%������Ƅ�X�v���셹������c+B�~��ף��ALf�J�1�70���,)9�f���.���Հ