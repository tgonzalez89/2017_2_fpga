-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
yPVppnzh5QH50YPs+AoKP493/A7F+0fyb9j3ahyndBv2Y9gT4yCVJr28ABq1qiU7dTvJcM+4YR0z
uNmUDWzkX92r2ua7EYmgTHQ8EXZUYBXSmchCqLNm9K0G2F65aiaVeg/fEwCZfcLrSJ6wUo71U5J6
nB4g2Pv4XFIW2x6OU8gQal0K435vdMKKx9OKVpgvFYIYPY0aX63SZ23ZYKS8/E0CO4hwxwL6puL1
I6sWxweoRjrH050npdwhj4cK6GDxoyp8oinUipKh8fEFr6+yEgPMXi2K85X0oz/c+1lKrHFGbtWU
791qZ3qTX2gxqlVI9etQYUg/iPrMy50M/2wclA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3632)
`protect data_block
WCYdIhxk36TfvtSpjbqe+R8xAZqKPicvfwOLNDzmFJwuXheLuZiaTs5kfay1Bo1XunlXm6tlB8Rj
3ZniRthJy/Vbgh9E7gq1UQKaFgvGlB2lk6GuyjhaMNpBnZD8oT955SpEtC+/ZVnV1AgMud0DE0zz
aH6eLIkm9uOanHLOzTl7MKxD1SVVCmBPHqJn/BjNV6m+x+XF1OXGsZ6KUmvoZOAwBPKsf68LB3wb
sIrKgvaWlStF5AS4Gaq6LxC68ljbxj26HZGbKfmG8PR4T0HYoNcR2qixzeJ8I81M2IUSmRfA6jox
J1NFLnkc+TX068eL8VDmBhxJ+AtAp53tlUulGlEvQRkMQiEN7++neCH8dlr0Ye5KHy66ZO6aY4WE
rY+Njd5BMkcDj527ApM35sCGTLKtEa952BtmntvNuP8e0tqkA9hVv1bqJrgaIR/PgeH/zRVBdolX
JJkPuFobpACgOI4Ec2FI9sUwhT/EYLqImfnzLYasC4ygFPnmjvGN+LTXjd0AiIu3ulJeigy5sk9J
+4cqeW7SsfG4+jGdANCldFXamSRDciNlMYFtqCVOvlEg8y2jo37Ky/fSMIOfKGt9c2lcdlgTjskf
OCuksVFS6x25o2b05hJPCLGUAsKkZrWtH7NQHEjVdwm061E7YsvPzz/1RFnqtrtmMqUJ1vtRpMmz
CZCFrODmcs9OSmmHC86M5qe1HV4HFLYQ9KCgcIyxf5cvhFS4P5LmaGVit82rx9LTtLSW6VS/mkYB
0oY0GCFKP56lmkhji2clWwjWMNJQykuhty0HPNXMYKbXIvhaLm00m7dKJE1lNS0zizzx4t9RlgFu
vJOt5oszjcS/+0UBCIawSN46wNWohK6V8wNqy3K/VL9vgeui9qZ5y47Un/zQpQrbJBa3/GLfCTQf
usjpEGJp8T9SAkNsUr0YmOr2UJPs6GO3s8HlYhtQdAJpOCXQIWoTYTsiqgGdm54ILWRrX0Yeg7A8
UnTRUY9AqMTFuO78AGVoKE/lzCq78d1sYAmdC+Uh88+QFaoSuybky9BNEA8Cj8pjCb877ToxqFWd
QTtjEBZ33FrRgDisxHUgOq70W0Z60JM6lLjKXAjU1KP4By+AnDAEmEY2sZXgFWG8KZ9cRVASO8+W
5lqUBg60Df7sHuE/27JNDVntWNFMwSVnWnqr9ubl1cKF1w5dlcpwKtY3CTuGJR97myJxP9INT0OF
DiuQAUI+zL+S3uTlkJHyD5b9JEchof6XSQh+XA64zZhVzIr+5z0lZhh5AoESqlNgaZ2UOOKHEUxy
WPSQRxxCr2IEz20Gzy+EMGjO5DpvgQBMx453+jYOsxvjbF8/dpiXHSZKg/9AHl0fXsqqRHqDUnEX
jDchV/GRcHjXc8RF9z4Zs+y1Cdu3CWnW75XPiJHz/YzkMYs29VPRGOGCxLqAI/Pav39+zCFFzTaa
Tihsh6nPuDlTEmxJSD9JpFR9QdHvgFfFWB/Be6CF8eOHP6j4MrlW379VN4oPUyfiIlSvIMZdJtfi
lbmN9qKp6wiPtFy2LDcLye1lTC9ksdZi2pAARySdxo5KIWSminrbIhDGoFjfqo22RP3FxrFI4k2X
c0IOEFxwcFnkdsJB4VXAdWotncnkAUnTeytKFtT0U7Hu8N3CpyJNso/iRCxEYbj//HelZLizbJog
7cwzYuShJG8WgHmLJNKlCuhFcb+glIQe/cLnArcGUE+bCJfYxzXSIoAwn7iFdT4F91b7MpZdoSi8
NaI6h+aax22Ds8Gq5pkg1cZ7EpgtCvmv9DNAhcpJFZFfZm98J9s0tUmMpjsJWbvTLXorctiREV3A
jc/SK6JVq2rYdChmyj/rv6t8OZF+OyYU1HdSPhH9ihD8cx7xXFrrd9bXDI169O2ByCtjQotkFfDq
9c9lsY5xXl9qm0C9fYGdpPX5DsXAg4odYt1nP3sh6xdEacFwVlZOHKlb30U4VJ7nHUoLjSUOq6p6
UueY//yM8s2tpkMxpbjZWT64qXgj85au/Vs4Tk2l+NHa++O2lnSxt69St76hFzG08v5pvgKvW61v
9wssveGAgFytGOUGRtIPrLgBUs2R7enIgF0xRij7wIoyqiUbtVPAhRV+fo5mLQ8kcF/Sv03xZfsW
M/fpAU+PPuK2/dsd5KqCOlQJtlBVTgOi/tkDM9A3IgqlmvPmg5jMyP0lmMAljf5QrmNfTId7E5W+
3DoJuynC1Zk+lkxZVSL5ZT8YmQOhZFtSrRwgeukkyJ3PcUaRh+vgY8vLrUieMw1RgC+sp2lMYKKE
kEuMOIgdwUf8X+ji6S6rg0udkQxPvkGS9e9bjWHM4N3eTN9b0cCbzGEetJnIasjf42sriIfsR9Ei
k06ZCdXtj8vll+ZkvqBhwBsuRvXxAoF+rUaFX7W3cG3pRcmNU5w/cHTBlz+6S0uE8sY6B3i6w6F7
yTGL8bjhY3FGisJ+oYm7jNMVYIaqvCT+WR9hS50/vemGwNIlVGp+DQzZMM6KtX74sA2eup/Pv1mn
tXW62Mrih9Eemqwqh3UQzmPBGuJgohXlJqsBF8JflVDTJyBxs+VIyriIUOVdZLCcoR/1K33W3OjE
AiGOQohrujdIlV2jdLqcA3aFXQoaIRSoPlM1HQu8ONtk+WxNK0VOXW2qLYexDzo1DSU9oOMaqGGM
DK1c0O9oq5nAqHd2J2XB+PKAFqaMgPO2RPSCe2E1x6Q9s729xK4MaJp82NRX9xpducXjIcsXyeP5
YxpNWFnAv2Ptco11t4hdwEIIkoomQjDSULMVj2xL+RMBIpQeylEwROmgS9p+FqIfW7FBOg25Omz4
4sgVhLN/YsSEE1FeqrC80C/uKx9Za0V5F2QZa4ZQrsVPz3AhcJ3jg600rZ1i6eYqfb1U0oX8xmSL
4sQHSQsZt0yrqxA9WeqCtxZ9lxEIU+7Cr5CPXZctwC+XmuJ1TahpFkOFL8OOOSBQZsRBFL6t1Kgx
VurClJifaEc1hgfWeFW5Ufo19pom5gnbd6Mrz1H32LanlHgTKXYYYYEPbJ0N8P744+4KRZC5rmeH
2eF2MO+SNLkoXUrHMK0I7QaMGnJVGlkDGxIGb1ZiHk3GyuCTKHYn/gnOmRqwo4mpdYB7PpAWYf68
gQaq2PhJ1JWzrwU1MTWxoidbyEjweZFcTr0VwenTV2MsNWPgCf7ZuVBt5hYYjQLEw8Z5gLb55+Ha
S3KwmYJ7p/KZLqZdIyo6kZOoPGKSCAwNu4SMN7ZcZx7vuNm32quOVjYPdF+HrrlOVFqLKm5qhG1y
W0foynXSEKHyWgp/K9g0gauPdfIZL4YNDrOcyIW0qdb/9IevevIp4LqbEuh4hzgzb6RpIby2+1FY
Y6ozKvfuFGOGyn7JFGJGSoqKPgV7lZcFDHo7wBABo91JBtRKjI5iihq09JEg2EgH8mhKQp7YA4SB
Q4LRxc4M6sybxmx1t0jOpPlksrPxFiUZ2awecsfmtQtEgT47VaKyly349lGqC18zqkApDdjc+xcy
QEiQp0LsQC2X1YIMm3DK1N1XLpgOtZ02JljPP7C3vUClkZm0e3Co81q3ka/luHSAgZw43nwBywrg
/3TZleR33GRN5oB1d2axEuOlhMxQa7eghqYaT+qTgAttIalsgwhCjlZApJQQoNF7YxrXg4YJXqtW
iHWKVVTHaMFbWqwrgjswFxI4Qe0+Vh8zgdKzfXmA1RxMF7TaldCl4+8GvsUMe+zeoMIx3iQ63Xzm
7Mpt+n48KUu8rDSk4T1rZcOeGxlRvY66gTWVouy0bCgxBQtRnSomPSFMamEOddbT3FMk14EWtMiN
TwutklX0i/0e0YouFnW2UZ38SEq8pd5wicrAmOWaRru4cuB/mLymwJTKd0z1HSvLw+ILoiF9ZUIl
pq76n/AmfL2NHgPWhD1ghpf54pMAwdeaz7qgzod4lWc1fEWRXTTeG9nGUMCxq0ZLFF2/O4mdvXZS
xXShzlmV3HWAW1nyU5HCFYyIYTybXg/Die78FWOL9GvLObfbd2opuVpFZ7vdqh4RkqkRoUmSVBqa
dfX+79XNtGDJIi0OHYN/5MBSNrAV3/hfd0immChp75VV/WL4qdc6At7Jjy/jKRAR3+hRQIsbL+JJ
nM0nlDk7pkOsE22tqwwgj3tY2ecu+45zrjYoA5yl1DZN/I+cMxH1vtU6umvq+pAtiRUWy2FHm1JD
ychP3JlXpYD5908FF7UV4gzkMnC8U/G8gSndI3rgLjOFoQvpIMppgf3W/bICqzLr2hLIMEpZWwFS
NbsRTqbc8YX8Dpen8aZ1ZuvwpMaqDC6T628ZHJF5SfqLI8C5lCnt7WmsMI4Qpz6n7FrM5xVtc3W/
vI9Nf9kcvWMReo9qB9mzxbytDzm/svyBcGy0V/CjuGNCw9GnL8GIQjv3KQILoAYCEG9QCkNzB/Th
lTFQiENT2qRAHEJiRA/thqk7aohS9MSoYF6mlSIamS6gkEn+upN/LbnZ7X5RNzXlHBUhymc7YiRH
utXALyVcLZ8yFRAvGk7w0czikKnpW2JoDLCdaH9k2Z/Aq+gROrrIaYmacg5N3G/HrJ1ld4Fu8Ze/
PJcaTHRgB5iS8DLjjdoTJ5/htZt1Xpac5uLihOAyMbb54J6TXmQa+plA1wRD2hnA+fnVbGfEnZwH
DSce3j6CbmQhK5STz4PkCXCGkp29QoW22Ajb/svUJPdr69IUpZduKSGQtEzPo8Lzf57coM3t2AxY
RxrP4IAT7+dKfrywQ+ozEY1wF4irz4xfCl3XQ4tCH0jGinn3yfWYsFI+wOCwVbiJ5PN7yyOWP0dt
nslVNgbPQGeKb7A5AxumCtdBOBcMNyv3aAbZ/aFR52HfY9MsOzNbHlU=
`protect end_protected
