��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR���[{�T���CK��TC,���:�
&��d!��]9�'D`�"9 S%�aQ�`!�6������V�W�l�a锦E(�\gC�slu�4U5=1�N�m��l�9ў��P���B�@+yg��=�}|֦���ָJ��^3^|�9�嚯�� G,H�^>iw��xnE���zЫ���8r���0���|�,&��<!���`����ܾ�z;M�PL�f�Q�!��6��Dl.������?�v�����W��^�M����@՚W�����h��L��y�;Ґk�`� 	��ϩ��L12f��h��;AP�� 4�`��]I�Zsq�)��b&M��&��8��C�-n5[�HW���!Z�Hc\�X�t�r�����޴9�:��.��]���e5e��{h %A�!ށת�M��S6�m@k�E��G ��O�=l����٬W����ī��.֎:�ɿi����¸^�E	�q|]�z͝�����"Uʨ�G0� �8��Q�pw����)81#7A���){�m��i'�#"q����x�XvF�˟&-�8�+yM�V�����L���q��.�A|�-u��Gߣ�����3�POǛF���#��c`:�Mc3舻V.�3z�Ww��e����𦦌>k�U��q���9�v�H���|-R3t6��M/,f�C����%O����"�Q@!&�:�AvM�f�*��ɺ���e�5#��3CP�h���&������Ł���wyϒNN�m������>�c//��pV5~r}�ޕ@"�vC_��ߎ'�����_r�f��Tro����T�Y�z0Ι�x�=]vޅ' �Ic��עO�]���`v��8������#kV��@������1��R �ĕ����!��̘Ur�s��f��~�,f�aD�����al���cP!�Fz�.i��~C��[0�9��u�N�����_tkdZ3�W��X����$���^I;�%� �����e�º��`@�5~�|nǗ���ú�[�ף�wA*��y�j���i���ԥ����te�}�u@W؟�J��Z5/_
G ����C45�ߣSG�V��pZ�ؐ�%�|~������7�hgl�F�`���Ë��=*��Nн�ЃP(~v��%�f�f�� �� MC�t;��>D��n���L ��ˈ�u���xQ���='���{�!�|{�SzN�����lD�n��)Q24������< �f_.
�%�"�$�k�9�.����cg�D���	?U��c{��ʼ��!���=�;USY���M�і�����3lЏ�4���^���������I���;!؇?�uS�BPD�^H0q!�SU5��$mJR0<���=�=˴�A.�־�6�+`K)t�ȋH���YN�O|��L�䄼Ќ�Z�K���%�Z����t@/�T�����z�:�*!�:5.��l�"�1UHM׫~V�B�/}l�h*·f�sgN��Ғ�B{�z�wO�Ӧ�*L;�(=��O#Sx�o�
^Y����#��}o�O,��P�>W�6Y�l7W����t����^[yB)�V�mؿ����-X�.��x\#6�����ҥİ��e ��]�P�L�[��կ�����6�cA9�˞��$�|�=�ؐ���M��MJ7�������0b�QR�B�~$�$A�r��b�4n�J��^t��(���^����͑����2�����Z��k �ЗR+Y�1v;�/Ꝋ�2Â&*��K�u�v[�u(�s����G}uol_F� ��
�a΃nl�Nr/�9�Y��5�n���#��.u�ns!����Ls�g���6�����h����5���'��~%U������]&���"8�M����/��I�;*QTZ`_bU��ݘ�x-���U�-�M���d��E�;$]��a�M������sX�����zp� �U�c�/�e#�#�p&���>~�r�}Ge��ή �0F���8&l4����kۛʿzۆ�ʩ�������sVV�v��	L�}l�>Huؑ����v�� ����q�"�;:�K�������!(�
=42Y�sg������^7��<���{�,�g��W�`�ț��B�#>D� ��縝m���M�Yr�R��*1/V2.�{`\�P�z����N�iX^|�3o�����3v?���M�S��LZL�ܢ��6�TJT	��I�,�!��^��>o�F�*�?t���:B}�[��;={���.Kd�oh�?��qPt�zDqX^����79��jc���������g��&W���k�����vn2T%�y����䛈,v�����Vf<!�)n�<+q������,BC��������� 4gq)t�����o� �pn 7ff��=��/�MĖzӒ�-�5"�wFù����qG�<
��Lv8�̰��tZ|2f;�sY������n�H3��?5B��0$l�DPH���|�e���7�F�T��7�۵�(�<��$ߐC�Yg}P,]�j,�ɨ4�\��"�H�<���N��FO'�'�Iè���=��>���9��8�-� pYm<޵h��׽��)x����@o>��8íFR|� <���PN�O��G��]�	�+D��=�l困+�D^0�Y?��Ԋ�Ĺ�;�5oo2C�[וf��|˹TPt6QGm���qe��[m���|f� ��#Қ����Fj�0�����{ql2H�W���3{�53�8���xەX�j�i��r�фy��Iv��P��)�]�B,��0��u,�V8zxݗs���e�F5_�h�!�IuѹEY3]��z� ���D �	9?|�������Y�T�P�3���0��S'ã��i�Y�������8�8�&�zR�u��I�3'������L���>uD0�.s�g�	�XI�2�������nf/�ޝ�k���-��/��:�F̶1�J�zܜ�ǘ&��4Ӯ�lN�9�'Ľh���Y	��c�1V�b�D�<^�'��'K��Rl��(����O����ů��|�i�_Vm�7?���K0Mɷ���1N�����������hK��_��k�����> ��
�'�^3���yO���P�A�bԂ_�-z�lٛ魉L���PLU�Vnh���0��:����X�^�U�Y;�k0���aυ��:"�D�!�c����D����Ai�S��@��`�m������A�h iy-h��_�	���]���m"˝�r�D(��L��o8��DxÙyf�__�NQ���e�Wc�%���{
�(�mJ�]We�C�N�8(N��7OAZ�#�(����Mó�bȲQ*�r��s�����_�&����[��>�K�:��0_��a�S���m4]/�D�}Xf��縕���}`�� �U�]s'�3v5� �#~��v!�ٛ��]�p��;ŢʅS���
�/�"�>�%y�Q���/e��z�^2�+�.�Y��`l`����P��*��Nw.p6�_{��<IU�ӋC�`X�R�yE9���`]��q���f��n��3;�K3�7��c'�C/3+�&*M�I88#����:j�u?����ŕ���&�[��̶vZ�P���E�sH���x�b��B׾����j��s����e��g��O��'��J]��}�{N�>^�pNN����0��*۞���'�(���*�q`[z��iT����$D���Y���5����u2��=0o��P։�w)��_����qaқ����A�ӎ�����Z��[jL�Sʇ�)n D� ��2@c�ٙ���T��h�	^��47Q½��p�5m+6�qX`�S��B9�o�y��YC �2o8�w�K���'1%r+��������QJ&�䍸}(Ji�rؕ ��A(� ;�9(�Xw��)xmx��|A3?����L�@u�;?�;�C���³�/\g��.�Ns�xq)u����eԯh���"�0�=+#�s@�4n7O�E����{�q�\P�r�p�h:D��(B���L�lUE:�4Z<k�*�Cq����$/�q:�Ʋ���2Q+yk�A�w[���0�ǧ;�t�n	���=R�h��Wl�2ڿ����[R��q�V�=���>-��,#�D%����_$�!�V�v'd�SC>���<d��^����/G��yoׂ�[�4ڸX��W@���-���Ԃ^}-��v��-�e�����Ә���>�&����o�g1�Y�2�nd8a|P�g��>$oF+����sՍ�_�؀��q9�b��B�Tu�N!V�!���?u��T�(�z_D%�)����ƍ����e6MM�����O9�c�z��:�S{�	�%�;&#I�>�����C#�S���1$g;��DY���g�=�3N�O`��A�K~x-�FU��a�y9�	�5���$>�tyC��`���ŜS������j���~g�Z���|�eA][���i�ңD@�+,, �\��6 �A��1\^z�K�2�����JKU��@�@Ḯ���Xu�)9�m��xKmz�Q�+��<�����j>�|�2,�n����+��o���j�aaŁ�MY�i�t��ϕ��L�aXe55=�1pl�k�͕�n^��W�6�,_בbV�i�]�:�O}y!v�4�3 �wb�VA*�B�G����~o�Y4����3�G��+S�����4� U���'8g9��h��O���6F�F$(�d��F.�Z��lu濔'�T�m�^K�
_S��h*T� 2��,�\��.$��w\���X���"_n�0����K� Y�@�M���},@�x�0j���>��K�m9l����D�J�� �:I�p��	�S��}V绋����(ڙ�Xzfn ��(��y�NPlD��\�m����U��b4;g�Iw�T[n\^��UP��[��{���@�8$вrI�p�G��k�Hx��:orx��]c6�4��棬8�����Xwo:o�K��I��"fY�	em�Uv��F����@�����Q<6��-��4��e,��ֈ��,%C?O��M��.N����H8q6�c���M�Y�zχ����Ȳdn"�gᩲ�|Tb(�d����=�a'
7�1����#=��g��.P��R��I#j�9���}��&���MH���y&��m��.��t3��!d��GW�k�Y�L.]���F����bW��n}e벱���࢏UG����(���Tו%�nR�=����lכ��4��k�����-��]9�3�Oce�p��\ц�rj�-]����R�Hv��Mg�d>��t�Z9J?I��됰	1*�������ݻ��q?v���n�0�9�!H�c�	�i]8���C�����o�\{�T�W�1����~eDF��)�	(B��3_��ؤ��<�sF�9)(��~��獚%���h��!�(�T�9�����,-'���;N��/XW��!Ǵ����8����Nǘ~���$g>�ƀ��}v��hÞP�g�������X�`&��:��j�LF��cp����ЬC�eh^1� �W����"��P�c�½�rG�$�ܤ�_hC����
@z5 �t�'!M
��~ę~���O�z��Kk���%��8ڰ����u�A�|h�hRHf�{�ǜ�/��R� ��y���]~u�>���j>�Ǘ�1}4��LL1����Z�+Gu��߾�`���3ʤN���Z�T�M�ey�Iq+�^���4U[�OP�9��Z��.a}S���z"Ɉ��F78��/����X���x��A&Sį'�۟�"��"I�M"���r-Sb�ֈ�c�6i�<���K|�ӑ�|�l���b��E|V�Ĭ �ˁ/'��uL�k��\����Tܐ���wDy_�j��K4�q�-A0w��3�a�=gV}��j02���+g�1Sާ�����}�X^ݫ��+�L�pe�Z�omE��d�"���5&9*��}�9��`o������*S��>~&�!�x�1���ңhl��-��o�QR��/�)i��E��S�B�vЭ��p��<����
�D���1$$^0߿H�b1�z�ᒺ�������m� ���R���k���7^a$J6���~�I������˅ȖB�C9�̦	c����>r۽��;���-~c0��D�5�OX���w/^Dp����NG�ݦ��7Ii<0��#�rU��7?�#&>�9/��g����Gc6��u^���/�^�oZr��������P1۾}EZ��Н����ٔ�?u���e���d�͇��0�0U�p��_7�i�[�}�7����TziN�9����m�����P�	����	�l�j��rO��л�vo���$�K���i�ȠB�a��$�:M�7z��f�s�b�@��,�=�/L��?�&�l�*l�y���u��);�Ĺ���\�f��H20���C�,�4z�����ҹ�
�k�N	�7�k������w̏�d]S��%��5�`r�ir�W>�{���R��֌DE�q#�<�nrh��Q.���*�sTy4:E����;]X��y�#a�Zn��7�elX�{2�8esgE�~��y=�����\���ޒ���hUt@��D~�7℈^ɞd���K>`W����Č2�a�H��"5��7|/� N���1���S.�?���쑅U����4�T�;٠׆#��P�iM��O9������RmxD����1Q�,/����0����p��R����7�\|X�$�di�����
�h0zη�~̬��{��֦��>F��Ƴ��*�@�,'�$�>^��1!�3Y���|�e��!���M἟;�}�O!<u�jw�hn�5���w�7��)]2.K�\�Y����`21硞�Y�`ᴼ��Z93�2��±l|&Q\#Y�m���5��\qoF"Ԋ^ ����:��k��T�������s��V|ZO�7�Q(�j�tZ����t'FW��Z��A17W4��$����(I�6��6v���yO5�6��\�k:�z��4�4)\�8��C�u�f|t�Vb���d3R����K����?��}���9ݍ~�)`�Nq�B��5 
,2����a�NhC}�PYJ���^���B��ou&��E��w�t�6��������cl�n�������¡�*�gd�G*��0`�����w?��	�J�:*H%�	��4'�5h�7�؇l�aCs�9�Ōv����3d E�l7�UB8��`�V�U!�#8�J��E�˂��I4�g��]���O�4f-�'X�7��ȷ ���NMO�il�-��'��U�+�G���晎'-��ક�sǷ�e��Ga8����⚺H�M�8����ݵ��w'X��<�I�����o6ÍP�9��rM���H�K1ku)Ꮿw"F
�iI�O���s����fI��Ď��D�q	�2�c�Y��[GV�T閖U�u�Ԯ��X4���ޔ�.�i�<��XϴѺ8I1����y*6MȨ�vu'��JS�Z�.�<�����\���Q2Ŗ�yPj��M<�~P<`U�U.���U������}�ʞ},c<*hkt�q�_)8^A-��R�{��2ڮ�z���ڑ�!��d��\�C���5�����ˍt����]��6oȩ�OH�A���Jv5�p��&��ކ�;�R�����¸�P���noi5پΈ�_T��x�<$�>q+(��
�彙��G8�p�&���a�}+��a._/(�z3�d��ܸ�+<�(ِ>��P/Y�5F��%�Ѭ�5�F��<����ӫ".��U��� �
ۅc��"S;i����>�>�!����Z�����Q�c��X��p���%xѢ-���j���HMџi榽��$��ϗ3b���9���"!(����Ddu���Bl��`-Ȉ��H�4��2�Q�V��|��x6��"�I����)�YT�a�9�)�hY�;�����C���r�BMsڬ;^�)5�D����qwܡO<���ޑh�����z��Mt͎m��S�ت�U{�Q���u@	l�Ȉ�k�L�x(�zN�kR��4���z4C�#���z�ȏr���*�>� ��֪�����h·��ūX����D�Z\$���<��7Ul��� 8��Q��l�$���z�n>�<͉ʂ�6�΀����u[ţ����wTu}�vmƑn�7'���%��#}��g������G 5��" �@�{�ǠzKذ�Ҧ��	���G��`��*���z��?�����xH�pC&��f�yx��0�zfu�y�}vv�}�eQ��M!唈� �굿�j7O����'��ն���@�h����,�-�38��[E#6?�@��I��`a�]���k�$��~r��)�UA�`a��xml_zx�V`B Xb���u}��k��p�� l�} �PZ����jꀇ�7=��Fs�W��|<.�W.�T�#Z��z�Ջ�s�C�]7u֜��o���P�r�6&3Ɲ��.˵|��b�p^��~����U����W�������ڊũ�Z��h|ƅ�� ��D���� � *N�I�/����Ϲ�� ���?.5�0v��x,o� ��j#���1r��Ms���u1HH���&�'[Yh�蕠bt��q�o.{tpۼz�X�̡���ߨ,�2�m��gq�g%#�b�~JaR�OT'⛘+��3`��8�"d���� �QpL���U(QM5�����ѯ�L�qâu�5�]JH��~u#H9�'�&�㋩"寉�7d��U���
��iZݱ%&�HH	J�f ��WP������1��%]PQ�5������}91�Wg;�qcZ�l�#Q�+-�w�Ƿ�@/��!������RL�����S���[�)Wm/�N�l�櫋���(fɲ��I�r㦧s&_���z]Cք6����:7(An��ǾV�A�_q�$hۚ� �S� >ψ#��W�K?�B�x��2�qe|�(�P�G�x��D�Ǻ��&����C�}Eۘy�^�$��H�27nU�n9l��Z�w��d��!�Y�0'��k�#�k{6��avSr=���#���$+�X5���S�)��i8M��|>�vs��2��Tf�{fN�L3��<�ڢ�SM-R�'l�8���ݽ5VJ�q��՛�l���,��V��[��PE���#Y�m�*��&�F_��zu��FR�(@.�P���!58�:{t5&٧��]箤�V�\�sK�fjp�B�~�)Q��t|��{��G�$:jcaS��� Q-�|,/��J�S�XХ�D�2��r����W4�Z��X�ڞ_{E�yv��j)"�e7i[��%L�#�.�g��q�O�y��'�(3�����M�@P	uF#Tkm@~	�@��9s�k)���Z�G#�F�P�r$�]a���.�dݧ/�^�M�g朱?�)�����u��d�\����(�ܜ����a��"�G�VB�]Ĭ��:�ym�D����w1qd�N�\I"+@Ϊ.��Bu�Y<`Z��,�!p�hj�S�	j����ߞ}�s�Ϲȍ�R��ώm��E��,�ia���pk^�wm{�#�WYz�0�D��^0�*.J����R�r���q��!�Q$��f�x���A,��I�NH�.f�������p���.h�������s�=l�;	7��0�t�QP���xHQ�.����"Ë%��=���p[��(	?L�љSOm�˪k>;n��0;���.�x�L+c���(���="�݁q7�1,/�$�����g�P����_�b(e`a��z�=��zl>�K�:B�G���X���ʺ[�/�Փ�o��O�F:�L�Y-Q&�K���]v��ʙ��&�̸�dᘙw���%�ʗUunÝV(�YLK��͸��QJޒ�G��r��P�/�s�3V�Z���y��j?ꉍ��X���|g	�"�vX�u�&��.��@��ύ�㉄ɍ����J9@M��ҏ<lyr/*��Ʌ����K��3�� B�d"s���^�ֹW}��G�إ�Mr�|�Ÿ-�G]0���;Ӄ�>�]ʯ���p���Ϗ$Y�#m���d_6�����\1L�f=斳O/�8�o^���Gr�Lڃ�R�@ꉈ4���-\�	��	��5�q��7~�I���H�DLn�9�ɵȥO=J}s8l!W�Y3��u�yB��& !����	6x�w��KPS� ט'��#��O5���I�[�1�����wOb��`�H�u�[��Ŏ�� ���0��WU�B�˹�=/l#kԷm�O�Z���1��}��*�,jq-!-�V��q�!��f#��|_��-�{�uO,�'�
���1Nv�Y�I��n�d���Q����z�����3��G�#T��A:���Bb��)r|ɥ� c�JH*��j4����yb'����&<�v�`\��P��}�vx��?��aE6$���n�O�[�� ��,��4p��R��f{����Z��UZ��alLe��n�}��wJ�g�4J����
��}���J��)�BT ꋪ�UG=/�<�5eî�p�[��Z�sN�
��N)�TnP����B�S�L&,@p`*I7d��A��J�^
i���t�:*芋7[4��7S<��B4��Y%2e>�vA��I��:m��T>�����N�Ϊ���1tx���o����k��xĝ�+�'���"�����Ee�_
ZӰ$%�;WjO���!��2���<��F{I�V�K���zY�	������u�?�2����ZS
sOYe%���@��ȵ�q��hN�rnX/޲��M���*��l���t9��y֔�#�5�m�B���Zh�Zv:66Z�o++Z�^�����-�Hd�-:`dcPak�[�8�G)��Q�#�Y����D!kK�����kJA�p��9|���"���Z|[��9�~�Ko��f�g�Y��o��m��8���3U���v!
 �T�<���=L��OT;C8*J�TB����m\��<��k�6�9{)���[b�Y���*����=��&�eD��,�]��z����W�����lt�Q�?i�k�{��M�B|<��P9ȳ�I��s>���Aa�N�[ⅿ��4@^H{hl���
�cBIעK�ǻ�� ����Dr\̠E5M;����Բ��b�^
dn,�qJ�6�N��s���=/PA�M�4?B��N��P��6_��f� ���XFʹC\mc����Mڜu.���Q��K���ʩ���H�`<G�ۿ��_2��d'L�:30�$ypv��-}9|癠.�6�8�7��:	�U��4V�MQk�}�1��L *nbO��x)t�MY���v��+DF
7�6{}-���ɫΖ��蜵[���5_���j�>W,S)-G��j��A��e�g��Jv����W���5��z^�"���+�V�B�ˮ��̗���w�HR�45�����h<CA�	[�E�{1�<+�O^\��-Xۈ:�;!G��P��m����	���HA��p8�/�&�t[x�\UP�B#߹����aTi�;}h���j� �����c��1ˤ�U����F�S���J���
�+*v0��66�j7��2��)ZPy��^�Ͼ�AsI��e��N�F�D��?@͐U��6��
����ɻ����1��5{��C�:2w.�7^S�/.���{�g2�����.�I������Vӳ,4,�h
�0<�&-��Ż��J��bh(|��H
۶�NX�$V��Q;/Ǥze=c�巠�z��D'F�C��?Z�-zxT<�F���I�#;0b,�����!<���ΐ�@���|.�����k�-`�b[t@��M�A�}'i�����D2Y��������(�J��GV���>�������=�v1�����74%P�V��xq������VX�����Wz��O�`R�j�U�ti��[��-U��o[*��8�80�<0���q�:K

c rRY�)����fD�W;��nY+I����]nQ}��i����Iزā��T8yc�[����:en`Q�������=�w+��+��QZ�(]����CFB����[%���"^��LbH�1P?Z���G��(����}{H��x�l4�|�6^�Y���K�F5Qa�����F�K��8q�����B�V>�GD��ň�:۵+�.�@��˦�Ui����$��a=�X���{;Dufz<r��E���d�q�l���AV?N�JV��m	��Ӆ�yb8$|6���~Ծ�o�򚽯VCISu�*��o��LU�iWQ`��6B6�Hb����_��O����Ⱥ@"I� g�wf53���@��Ї��lH5�Mk��zT�M�t>��ׁX/+��;I����H�HY�%�Bh���e��� ��=~,O�o�=�&�S��^6绦�]yu��0'���=j�f�&T1M��/�,�������A+Чw��ph]e�W�
\Q?_�h�� (�s%R�z,O,^[�|ଃ�τ^�<c�g��ݪ� F���4$"3NH=��9t�%%A�J�u������"-��Mδ����*�-�5Yd��F������!9�^,�G�Ƌ&6��M,��.�����"�;���}�Iv`��S���msU��0�p�g9Q���|+݊m�vԠ�Ń���rek�dPȑc���ST(HR�b�%P���(��C��-����݈^�s�1��-R#���(�_k�[��"�=U�Њ�gfH�f��S� J�R���س�6�s�y&L�K�D�����7�pG����D���V�z��[W�F�c�{�6$tR}-SW���4YzRkFx]�:D�k�i��"�1��^c���W+��,��iFW�N.�*�i ]x�{W�c�rV�U��?~KV�Xwv��"O�6��v1�L �U�ml�u���l>B��	K���[��s�>�jߤ�W/O����xfТ�>���P���Q8�)�^���c�O��d��\Z�� �loη�	İ���i|�Q\Q�xxH'����5;M�`b
~Wb�3�� q�{����@�̑' �9�P�d_�"QR��h��lJ�A��=��	�j�(�� Z���M���?��1$��s�j$%*��A�]0o�����Ƥ�D��D�&/��.K��"���G��Z�)��U[�[���bla(�4�['�|�"��Xt��#<!��Z�*yi�qƹ���bB�0u1MX:9�5�<t����P���:j��r�DZ��V�R0,�g�Q�E�`Յ�aU�Ҧ�ki���&z]X8z�H/$D���9����u0`�U�h���������h۴ø���i��P��=�|��x ����~qa�$bf��j���\��(4'�c��/!Q�h��q�̡����ߢ7N�����'6��rڿ
�T�ܛ+}GL=�OpW�;�:=M�\�ѫ�}�[�jq��~pCo/U�r8�ݐSv0*�7��UtfXz�@m��S�̑%=����K:r�P����k-���esZ;SeG}G��MPb�9|N�p+�&��(tl�$ٹ�\Q�`S���܇��M�]t�
'�#֘�	�{h��TX+�|J�)����U���/c�\E8�V�DEKlN*Z1請@ny�(�2���`g橑�#����C���G���j��; �}�U���P)v��#~�&z`��Ll�
����s��k-��a���bu� �Q����8�>��fę���WIb�m��z� ����,���qmg{�w�x�����1�����d!����m�%��ZK̠�g�����i��jmnw��Β��ޥ�K��hc�J_q�!r�}�t�T���kP�M�V��g��%>�FX�"�k7I-o7p:漸�kr��]h�-�ˉb�{�1���FA#]�����(���p�l�H������&?h�
}Ȱ�Eӽ�Gd�4���,X����
�@�h��� �q�+�.��״�3 f�M�..]M!x@��M+
�Q#��f"�HI��H�E���qY׻�{���Ŕkz"l���y�յlE�.��p������,�	o��[Y����������#���)���2Vz� ��nB2J��D�R����Z����%˹�s�  �T-5oQL����kyh�ۃ���0z�S�2��^y�ǘ6��K������yN�5Up��E<ݼ�+�6N�Q{/�^H�(��[�����>�����bn��:�)���x�ƪr��t������v�z�TR��HJ>ø�Q�A�>1����AGUs�e������$�F"��տ'
��� �������e ���0xnc�.s��~�g�_��n��v|>�郞��9���H�/��d�'W��۪���]��Lo�L�o�OXa�X!4�gy�`M�Z�9�ۤ����YV�	��	L�����y��}�/��w]�ֺw�V�'���9��� �!�U�����g;�*PP��t^�-�0YV�||���m��% � j�{�7������f�$*2��&��g���y̝c!U$���q�Q��qZGn�5��@��:�Z�4�n0�3��P��!RKw*V�g�+�����&M!QGX[3�o�[����A�S�#������kPP7B�ܽ�Fa��j�9�I���n#y+(�N�C%�&�s�-���u�T,W�STs�-���>;��������CԼ������r.76a(:�X�V�(U�@����Y�M�Ē^$*�^�1vT�#C��3ԛ�.��+Y��+�-3AnG~Q�������ɹ_�z�略Z�$����ū@����K7O$rEJ���vm��׬>ʡ��P���as��N�
����d��#�Q�pz��N	�%M��9��*SL�K,��δ�ocL�#��T���p0��9���\�Nm7
DZ\�m���H$(¦-$�Ȩ�-}�P$��X|��U_Q9ًJg����qkW�gb��苘�fE,x�)�㍲b�N�
�ViO��8�ά>�Y��`���$^]�8
��gKWn1�D*�'6�?V1�g�(���z�_�l�v3��y����Z� ��aL����9ĸ������	�K�I��.s�j4]�K�"�8w���͓zgL�Vl�A�#K,�Z��o˗��T	S����c)����}Qus�iK-_&��A���,0�\���\��Z3��q�$��i�ɿnJ�tB��I���/��+t l���A�+��<�]�M�\��3��$��<Ci2�6\I$s�`��@�;R^x���8�i�+s���'b���E!4�:Ico���؊�$,T��Y�L������a3�z}���^w�%P��I���(�[���t�-2�	Y��K�Yc�
[�����̇�|�r��z9�J�Dg����T.�bY��J�uk;��bd����(�CɊخ>֗`
 ɚ�G�G1���Ra���G��5���W����{Ԉ�M5Y�D��V�8�Ƨ�i���6��Q�%0���2bU�/l��I���٧Ul�[%��-��?<1�Zm9��z�8�i�<�ۂ�-&���{�'X���IlIs��� F!���k堖^���񒹣W�_�'L)�#΢�;m ����!0�\5�7�S��o���gœ���e@ؼp�{�Pϥ�[��]Y	�W�iB��B�Fڷ�é�U�H�ӿ�c����n=W0�J�<eІ��z�TJ�R˸Su��}k/��Md��@�9bCx�ك��5�W	�hz��8Ӫ�Z��ʁ����hTxl��Q�XU9�E�4����$�P��\h����3��zQ�֜���I9֟k?WJ�p�oATS���OL���y��\�N�H&���X��W�7�A!�+�S.,�8Vj4�@��a������/�vQ�䘨/�cI�be��t9z���x�Sb�'��@g����w����j������It���GK�����x	����� �;�^<he�2�[xR��Q��;�w�؁��$̤�`���@�Z!z[��HN��H�J��<xҠ��P��i����b�!��DQ�n#*!��sL/Œ�W?d��ĳ�N��E!˃��un�n08D�?JTFSx���ُ�+�s���&�U����6b�_��0�%I�\�\rP�ї�h��hp��U)�n+���I��P|���*�s;�a-�dpt'T�4�R����~�zz���Ʊ��01���,�'bK�X�t�F��G�EP��s9����?�] �+$�ψ��	���`KO*!�3�����Eust:���&t��,�g�1j6��8���3*�S����(����&"�=we�<l���?b�fްx[_�@K[ۀ����K�>�Q��B��i�"-Lé�"�x}g}�ʈ�'zE$�*' 8ڏ��I��GѮz�>1�*Y�VY��~�xt��+�&�x���"S�!��%�Sq�KQ��:��B_���!�g�5�̕�jPT}f�- �	�Z.�y��}1��o �pdnuM�e���$[��D�7�>G�CPH��A�#�rS����.J��d9GϵحKl�����3���툓O67�>�rF:����������Bڰ�z
a���U&�s뗰=
�T�ET@֨�A��M��JcS�ˌN�CD%U�I�;�������kq���v1˄���2��=6��m��rp4âM`"��h��ZF8�>��N��.�����)�?^��iFӋ�l|���U��]_#L��t�I{�I��C}�����\ j��M4a?؎�HV_.�7�Ͱ�[^�ωļ�_\�Tn=�`��bo�J�i�t��ܹO�ca�5�I��5�J0��h	gR���X�bn���sY�<���-�y����8�nt�h?�>a C��3���E���޹t�9P�2�&46�{�.$s,�$�����t��'m�r��"��1Hf�ړ����0+��sA>�SP�TP���N�	���(c��a-,�����։լ�B�ȃ�@�qPI7O',�=)�
��g���H�j�{mpxM��:�oP}HQ�
�6a|.=�`ez;�9hn��k��CnB� �H��nF��{>f�/��RT��V�|���2)�{iH��Ӈ�Ǯgr8��o���ׅ�!�x�{7>Ez[A�	<o���������� 4HI���J��2�$��M^Z�z�ؓ����K����e�;�O�ժ�2_�s�=�����PX�x��01���?�����@�=�z��'�Z�[҅�0#���E�6U�����b��&ګ%D��0!��t������r�m�N
O{��4N�i��ς��3d�,���?V� ��$�ʚY-�D����[O1�\c})�"�b�����B��ӻ�U��קAJ�y��?TA��%|����AV���?x+u1g�e]|W�t������rs���$��K���V���Ɩ'��`�|Y{=_:^�fM4���h�{&�A�/�R|�XB���\���Q�ү��HP�Ev�n��^���l����{�{�c�X��!+Oa��)����T�������,Y]���5�� 2&d��8�*��Ȇ���[4�}���,xd��k��D���p�?u���{0ԇ���a��>�];u�5�`S�2��a.�8ʗ�'Hl��z�8�����l���Ҽ�1��^�!��=Ƿ7�@��ܟ�!�/r0%2Y����ɘ$aFЖ�����A_{G($Ԋ ��ʦ�*��(kW41���4�!��Z�m3��u,vp9�6�2��yc�H��	6/w�G��v�xt���#c��&X�� >�,��)G
�ud�qy��Ϻd:���ǒ�Kw81��=�Ƶ7��ۑ�:%GH�ʅ�l��3A0Dq�r/{,�ʈ'�p� k�`��3��
9���Ft���bN/c���)�!����.8�?���0�s���NH�m8"��v�5���l%��g!㲨ֹ�(�H�_�L�k��`��;��.���}{�r��K� � h�u��Ә�]�c�(���S��xq�&9�� y�oZt�Ca�6�=�z��wq�� �']0�6/tyʩ��
��'#�>�({�����n�i��Z���U�J�y*2E�-^�A)�ʌ�G��q��ó{>�(��8�R��W����S�z�iߒtw��Sm-��ɅK����Y,��[�ٹ�bV���Yf�KQV��$:��:+��)���[ӷ�p:�=|�� m��߂���o����R�+5�L�x��.t���00�p~��sN���@
�]"O�H�uA���cfw���I+>�";��|7re�zN-g�z���f-�h�?=�v-�8�@����I��)���8��%F>�J�^i+FT�l?H|,��O�'d5�Dsy��0��t$L�k�m��������gl��gtg����O�;Z=O���<!�e�tR#}P�����Z�������B��)i��@|�fDv����$Sտ�S�tH":m芷A5܊�8Wq�ݩ�w�ޭ)E��sX���/�����^C��p0<��l��.��!����֊�W�Y[&���E; Oo��A, �@A���w	Ͻ+��B��m�5�z��C`*�|$Fu�t��6�3+P�;�����[���|f�!%c{�f��6���rk��Ց��#����ٶN��������#�SvBu*�W9��v�0g�n�%	�%�o��v�����*���6���))(�}j0
\��/D�� ���S�w��/B���Su	u�/�6^���`y�GA�o���;-!S(Ĉle�֦5�D��Dp�a�#���~YAY���|�V�����-����m�H|x��5)|>8�#�.0d����=�X ��T��y��C� ��>Ȁ��Tt.>>
�����1͇9(Ӷ�<0\�&D��E{�v��}���C���v��F�`�=�������?aѳ�bq/��Xz�Hc�).UN2��tH.)s��t]vd���s�\�y��7z7M��cw^�E?�b���7�J{�5�Wcӭ{(K�ׇ�f��� CE���@���;��A/ǉМA�E��|=�ur���~����X˝��q�:]DP"��X����<p$e5����S;�ɒ�=�7��˼�X������N��ee;j;�i6]���i@I��豥��j�)��џ�@--I�G\��0GQ�Iy�D��=8�m��Q�_ :����3�Ѵ�8&W����X� H�|i6u�o^$�����v&��(K�~����|��^P	ūy�����{.��f
HaW,	?T־篟h�u�撤Mb��c';�B�ME�����v��x�	#�5�.�S�̿�df���~}��44X��W����P3)P��� "��nҿ'��*3����p&\<����������6�-	�%�]�ĘwiP��cٖ$�	� �o�c���F�T�H�|\ӍtE�vJ`_E��[d�-��g���J�d��F�G������m[⨻��%)����@�Ĩ:�䛼U"`�ȶ���RN�lO�$�9VW��MIX]�}F��cw�H-=G[������S�&36a9T"`�㾻:�H�6w{;]n,[�}�I�7�ʓ���4����W��꣖/�F���V.65�2���l��\�#�y��G
�$ү8ƅ�B�x�zq��"�앝�T���7KR���Wc�;�0�24J�lX�0#�AŦB��DF]�:�He��HEM�;���[`vp]\ �>ה&��H���r���aT��s�l��p�R��C�G�%���N���}6{�]hz��B�!�2B�#Xrd��7�LKO�6��F������	��m��./m0�@��r�1��u[B���H?�0.p�Y��R>n�L0��k4�¥5�KD����)DO�	mY���g���[|�����gv��Q����u�Р��1b灐�Al�>�=����׷i�|Q�(��`���5��'y��N�7T��hJ�1�uN�P�!��/���!��?��ap *����S�{3(.��m��2M���=�A��;�W[z���h��C����O����Y'4��o�Il<�j����,:	1�Z�ܲ��ܔ��쌥(���P�)�a������@٧�z^�m�c��>唉�k��tR+tz��ٛ���g����F�y��a!D��T�_�����GO����i��!�Df�s� �/�Ĥ��i4Ys�.�{R��8Ӥ�<�f���n|�w�T������^%gF�6Sb�(�T1��=6����m��bvc���*$��8���Q����2㗕zh�h�.�Dų�B��0Sۛ��+>��Z֮9�?����ɤB)Ψ���H�+h2�1Clq7C��~eŁ.r���4�|��:�䰄�v�i��"�g8�~�-����/�R�yr��`G���S�%�|DpUX�u7�XH��<��w6~��4�z��U%�y���iŖ18����J��V�TS����^��ky�����q�~Y��4�_���}�ΰ��Ek�~C�MKK�����aԏ��Ʒ�[j�Y) :���m���Ov3�8q�9����e^6�w�ۏt�z]�t�/�/����=��ܶ���� ͟��Vm�+97 ���Ɋ$'��%�]n=�!�ظ������#��	��6�6��V��@�xC�bϑ�K��Œ*z	w��f�Z�W�e�!^=�V	�L��˲[����d�h��#�Ľz�yrŵ'��`x �f��H���~�ƍJ��:��I�-����r�!K�-�R��Z��5vJ ۴0�lڭ/�qm$]!1����f���"qX{x[+��n�@$ hn��R&�ku���τ: �V|��pD9��=al�IDʨ�������T+r����ߔc��_E�B��H��� ?�A�LC�6�D�_�V��H���W�� d�V�!���e����^+\A#m�$�3��eT�����u	V�9oU��8Lt�9s�b06C�^���J�n���Y��P�Ba���,� ��pS���^(����� �k۠���9�.��,�%.)��
>���t�w5���ũ��'��Z�[�v���P^Z4(�s u���JǐL��^�X���W�B�vMUv	6:�v� �]��۾�s�x���d:��#�E�VQ��:��Am����UK ��z�Ӱm]]%�v���,a����˗�����|@!t���^�O*��f���R*���*y�����g��o�	�0��-�T>,c0���`|��Y�??AG�T��U�ۉ�q�n�V�Q�\�My�"q�m�C���+ų��{ M�R���y�k�%���-�M���O".���6Ln%G%��!�kDW/�o,��E3�/��G%섖��
�Ž��Z��;�Y���� hO`+$5�ט���}9�|�:4�w&�r���1��^�;�z����C��u���L��������iF���GlW��[�w��	X��>�!��΄
�U׫�g�|�a���7R�	/w'Wa�W�����/C�"<����Q�'���l��X��A�ԍ�m����WDl��o=��&���Oc���&ٟ��iә�;T��)�]h�ABb}�\�K+=�	��m����L����%��Y����.S�>��?E���l�G�HsH۔�d�H\��H�v&p�m���;���QX<~�"xO�ӓ7���ɡ	n��u�e���,���=�L+� ��5RL�=ԉs '������{��hM�ޛ������io�=��h�>g��z��P���2
T��_&�ZS70v�яt;�tt�$�X!e�#Y2'Z)�" ��:�gMyyĞ"s��c�Б��KY�#�4��7a�qT�|@��Cx��4�5ώl��{D����ʂF�}*�Pɶ@������lkXŖ�F��<CQ���c�
_��6�s�Ԁ�b�D���x(  pسM*A��>D��ͱDL6���4ST�`����P/6��i�=w�8��E�K5V��qI����#��v�p�_L����-aF�.��x��gH��y��p��P?����H�4��~a���X��O/�m�Z�\���BG_
t@��Q{+O�߼��H��k\]D�D��O��1��?mwU���,��5����_>c���Y˅�8k� �_��L�tW閫�:�������)�����]��(GL<�,���3��5PB�����0��[(�E?�5l�D�_;f>R���Dۈ��D����H�P
`O�A�2�a�<3O�J,A��7�Z�v�Ƴ$�"1/<Lb�ٷ��q��\��s�g�z��rـ�n�^v)L8իGFq4�3���N6U��tТY�o�nHE���SqrW�ݟ�bkY�Շ�(��+��J����7��v,�`y<�>u+��E|��.�`q�mg��P��j)���$� �p���?��{�oE����Co�"Z=�ec{B����O���s�s�p�ޣ%DW)]����T�Q�����pW�k���2̢O��/f�0��T�;E���*1�%�9�� &���!�,ꊙY(<D��R�E��?YR�]M�{16K (�xPwi�u�u�v�aֲT1_4e�rcno�D�2��]S	2KZ��i�� " E�i�G�N݈lǃ��u�|���Qdp�9/�4mj���?P V��k�mҫ���;��sj����G���w���b�� ��Yr2���ŀ6>���+�8�y�8�\N�8)7^,p����GoH���	�w�yq%����t���w�AM��D	�s���9�v
D��?tfW��ZQI�@�y]��]z&�D���)gϮ;�x}�YO���"u8��_��s�B���}�N$�/$u\4��UŹ���~���z��7�Э���6�#m$��W;
�yj�4�V�vE)�/�h�:�+��f�,�	�!���>�#.N�����#㪢�TA��^X�n�YPE�|L�%_u�M֑���H\<�y 5K����4����)�q~W���y�����Ȝ<�pi�F(���}�/�1KyT�~���U�D<�?�A+��7�J���↏���இ�2��.���J�R�Q�ޘ�J�'���$����$�J�%���ۋ2��?t��_.?m��Ƅ>�dfN�#f�0�Q��\C�\H~�(���n/�U�X T�S��Q�m;>����m����e/�D�1x	�r����,�f��$�Th`߸��Z�U�^��ߣ+.�f��i�`�/,�����.�U��Fxur��Ȇ~��4^�6�T���~�K�Fb0���0�"�F�Z�H%<���s��j��\eѭ`��(�
���c�7���DQM,M���Ӥg�놰�&w��Qi�\�ԏ?�(��ǲ;``���^�V1�Nڍj`8 ov,��k���	!�$tt�u�XJt�RDԒͻ�mI���g|�ͼC��|]4�Is�JL�A]��K�>�k!��� oC/I#�ٟz����$�Us̷v�g�s.�Np�	�Y��dZ�m�a��o�mO�Ǘ��"����A�i�ߧ#�)���w�O,�+��,�F�n�F
�#�÷f5�[���ʗE.7E�l���@���_Lp7��-
���S�'^��f|��JcF(��Ľ��6�;�UȁU7���*0��1 �W�G4���+3�*��x)������bY5�<z[���LC���bՕ��Ź���~�g�$�	�%vnĬ�[�w�����]�1(RL�Q��E��X��ݘd.�z���td�JN����8��R�I�.�`�>L����i�R'��q��\�!�	�Ҡ����ޚ�"#׭چ�!$-�o�������m髾F}B�Mz&!���9n���-�^�i�2�w�M-o���gu��
�pqhSR�.�hF%��b 篰�k����h��v�����-j����	;�L��f�c�³$Y[��@	K(�(�SvD�wB�P��_<X���a�&K-.����J�O2�ҧ,*�:x��
*M��ߕ�����r��T��Z�1v�B��S��Е���d����C���P��eΙ�m�RO�WS��8O��g��.w����t�@K��=�WB�A�0G�>���>�XR��)���~���ߩ�bts8� ��ddUL1mQȍ�n���+J��F7�טJ�CC�Kw��)�1ܗwNuD��ј]��bI�dގj��N�97�g��H�|�@k�^���.���_V����\�d�RȊv+���X�4TB�zO�!,s�g%��ʏg�~���P�K��`�J�Ca����Z��ţ[��4'��V��	#*RK�����h��!8	��1�ә����?X`]c�0��k��,�7Uai����������7wB-B5f|��w��Vd?Z�w��ai�$�$h���R�>��-nPC��;ʽQXA���6P8���	E������[����D�U����1����]3=s
;*�ͦ`�{�@�u�5?�A��̨|��^~w��E�2L����
LB�:۫͘O,��B��u�. ����p�T������}0��5��ܔu��yI�˘{�I���6ڞ.��-����_�ؚ`�3L�6n���h��A�9�v��J�>u�֯��zA.59T�@+���e�,�救P�&��3�I��%9z71O��5*�{��cO#�����n�sH����j�	�;g����{HV'��l�k��n�v*�GCG@&��� ��n��<�%B���X��m�~��l_1O�C����p'�6�Za�����A�)�����ous�U6��1J��$�}Cy��I{��H�g�p)�B���5�`����W�.M�f�%G���s�E�Z�'m�/����]�tYƉe"��R8�؂�<-w]k�#�3�(v�o�pUX�����^(�NT�5��x���|0���P��
�л�b1؉�=r�z4w�~�����;�H��������f$�P��2��sF�oI��}x��N�ǜ�/x�Ls�v� ^!�G��F[��tC۵��&n��w
1��]ĵj�3^��sw?����c�v?��6��VU]z�!j�g�y����N*#��uW��i���N�N�7��U�yD喸E�g���a;�zť�����0��;&����Oe�����$�U&�qY/j�Ʊ]ۈÚ3"�~��S�f��;.�=:`��i���j��X~�W��[�b����®c�������*~�){��P/(Y��T1�i|��/h�6P���:c�=�Ì;\�w�2J[��C%��rCP��FLx�B(F��9�D�*j�lW�el��vkSt�O#Mk]xݬȚX�I�u,O�n�r�9��,�����ſ���˸s��k����3mK�r�Qav'�lE
$�3T�Y�SD�.�&+�M�.6�Km�g��e����0���cs|��.o��AGjm
>PwC}`K��{�P���Y���W�_�D_۬�|>�!���h_���>M����TL$�@O�B�%�bHRn�ϭq��N��I�V|@Iq��Yل͌*�>< �<f�`�h,�ri7��e�K4���ǵf(�U�B�+�Y表�eeؗ�J��U��[��<��:[5��I/1|��d!��EQ=]Q�w�C�OE��^.�@�mW���r�D�)�|�q�_N��7(�yr�`@LF�g#3������{TCg:��^���=5�J��'St��!�%0�n{fGm[mf#�7��p7��_��6��:/��~�i��RRzgKuв����H!�����pf��Ӓ����{�i%�W��7.�����9{�mwlê�O���K(����ѧB����.-I����
� �kP:�[i�ċ�}Z�-G�\��`��C�OQ>#>�)ն��K]�ġS]��Jjb�[1+V|?�ǆ/r�k�tЂuǂ��G-zL���hjQ�Q�$70��Bu��l��S�/Q���؀��I5}�PT�0,�C���d��	�K�x�
��q��6E���1U��J�[ۨ���W�!G��ś�W	e��ͱڲ$��P0o��1Ƌ��Z�?J�v�9H�{o�2�y��J�J�S{%3x9coL_Y����Teh�D�C���q6g9�=>Ø(DqG���;*�FAbrO�o6��~!)|v�]x$���m�l�R�00c�\��>�s�֙-�Jj���?�e~1~.����cY]`4�UJ�A���C�?��7��߁��Iyա��ŉC��Ca�6�Q7p?̎'�Ъ�9$ªy��4���lۄH9��}�q�<|������uG)��m�G�G��[�|J*��I�]t₫�3�x�+mM	 `BVI��i[p��ƹ\�� �-��*�S��O=�T�~l^b������d�P����e��
���@e��X=J��%�$j;��`B����ټ�:�׆˷7���n��ϓB"\��r�A$�{�g�e�lQ䄪 ݓGA,1L1'�Ř�Ux��Y5�2X&�O3I��%[�~�:�[��!�:�;�o��U/�(N��Z�'К40�$�ۖ��5�S�`���S|P�U�� ����?ќ8�� �k2����{NX�[�� ���#���̬��[�X�;�f�$�܈B�B}x����Q�@U��f7ݙ�kzx�;�I��q��Z�ࡡ��T��Y2�Zt����;R�d��'���d\�΅�\51���-�T�ݷ����¥I ���q���,D6��s�ě*ܞ�}�ؤ�w�@�_�$2È�H|aT?	pMY_��"�yE����8���x={�6P.gA�fcƶ3�k��ԋx��c�si|(��+@P�Q����*��)��u�~)�XsB��W����bx=ӗ��\��ǉ��J(u�wv�k���Rn?����H"�&�n���dk����դ̖�0��$�|���s�D+����}W�8��[j�rh�������?6	K��|& %��ͣ-�e5`���r������RC��H���H�4�����XeŨMKiq#�٫�T~⁠��iG���OL �� R��4�ޏ��;w�΃ì���ѱI��i���M�G��E<ŊXB*1�hg8%�f��~�f��p$z���T��_˼�1�)RH�I�ԗ��xj:�v�#�Q�fw�,�l�ad�(����H��tI���"���P���\8T��,y����������S1IAX�AI�&��$��HN`�蓅K<$|�;�qxDT���@r��h<N�l%�� �gK��Fl�3ƕ��nc`��" ��)�C[Ҵ�\�(���>꯽r����4'�@M�U N��ќ�*�hۋ��ǹ��[�I}��Zt%z��8Q���*��I<�d^[���2)0g�H=�^K���'{l7�D\d�HhH6*ړvk�,.^�_7�Ի��h7ͤ!Go��k���� UB�;zP�����tx��7]I�"|��4=7£K]Q�Ƀ#d4�l9إ�D��Y���$��ƻ��^-Ӫ3�4�1E����,�)bB�Y�(�a5&���W��ڸ��P^��l5c��G��_^��r����+�ί�&�,�0}e�D����ygZ�E�kIG�k���p�x����d"��)�9�ʕ��G�Ow˧���k�(��Т����{��:9'\�Fc����lH�G4g9)�+�����L$l(��wfE��RH��俕@D�̦�Q�M1�u��{�������Ԙ��MY��Q��D�N�܉23XȇU[b�4~ޘW�2X���F�=C.�7k��سFg����VP��I��j��9�F���������<@��p(m��V��ܞ��}%/ |��um77��/J¹�̩���`C�7�]P�j6N,Ά�Ux�J�wԍʉ�$�ٍZg�=<__�O<�*�
��-cI$l�'}���k�ǲ��)%+�_���؀'�{�W�5-
����ú���	"����ʛ���ހ'd]1�68Hr�*�� ๽)ڻzY9b5병;߾G��r,q����O�Y���u�(�*+ �*fm�!��4�(�T�5���ݣ�8�D�_������]��7�Pɗ5��w�Q5��l�c��&!`��MU��p@z�4p�F
]iRjY����D���>�~�?V��G�
��,!���9N���j8�	��Lw�	���D���~:�q].�~@�i~�?�,��cXb��"Fc5�K�/��q���vH�T�v�!�V�9mn���:�C��laNTZ���wV��L�p+�%�����ɴ
���}�om�?�=|r���Á�d�SH>�	=/��H
q%��(����1D�Q��).�C����]`�oJ�(��g�����U��;��h�pjݖW6̫Tc�x�z>��A�!�Aqpz�C!�������Tv���3���*�X�u.bDh�S���rH�q5��aY���t%�Y��s�)�IZ�~=ޯ�v�-���;7iy�e�K�qn��9���	���4���?_�68��Q�-��8Hg�>�:o2��L%�{p��ΛE=P�~e�(� t�����)�����l��u�����]wB�=�Q�p�dL܉�쾕���#�s��MXrn���,�`���֔������}�[�.��E^A�W����^5�.��0�jhٴ]�Q�$�$���r����P��v�Ô�>�fK���g��/A� ��Y9�n�����/
 �aN,˾J8�4��B,�-�k���ʣt�/�8�d�����|
�de&P�������,�(Ur�(EP$QW���`q�ǛP)�����O�@��_?>1Ĳ�I�+H:D_��g��G5�u�R�������>�F�3|�(��l�PX����]��3�V�>��:!����:	���M�����������7;ȑ�n�ڻ����4��+%�)5q�"���b���,���T�Ms�l����,.��s'Y\{_�7A=�
�d��L¿u� E]��PW��y����#-����u�ܾ�@�����gv�[�θNL0<I����e!)�	��(k�!�3���`��f������*y+oZ��!�������O�l�b���,�t:���x1�]mdҀ��:���0g�H@t�`� V���'7/5M��r����ÌJ
�a�>�q �G;����1����,��$���<�<������+�x����RWr����*��Фʼ�N���!<�&x!�1]�n�g6-��N@U�銥���U�C��wuXe�)Ky�'�x(4����	��X�.#5��*?W��Zb�����䍗���A dc�]i�'�|�G���n�1����H��+�t�(ygj^-`�Uo-"��MF=�>���!�%�u�fZ��Z�	���2�>�O�sn�n�B4�R�P��������p��Z��̭�.lƵo�VGPmШ��o�W_ �hr᱖��v�~^B�0N�-�$3�t:Ԟc�/��E��Qk� V��y <��ŗ����W�"T�E��q��5N�����Fa�n��5�n�RB�Im�e/ ���%`�@�6�(�՚�1���a)���^!I5iO�H�s5�pt�,�n��!�E�,=]"�K�����_�q�JA��+����&�TԸ]�e�q�H��b�~��ϵ��9j?��3:=ku����j�����!�L�����y\��<����=�y��&���J��Y"0,+ٜX��z�7�rU/��2��f�+�ɟM�t��qi���Wqt�ل$*a}�e�fܢG��f���89?��5�(�D
Z��L4�~]�ǫ�m�<"��x�<t~_�w�.
�D�|BB��N���VYA����J�chG*�o��\�En���[�K�	��g��=o�O���
h�������Kj1�6~R�XHCw���F�ViP��|�z���k�py� a!�D�Ԡ�?�,)��x]�I�uӑ��R[��+"r�����¯�V��y���5f�R9�y�k���?*�K6-����"�l��p@�`75�C�輻A_=$��oJG��MLH��)"m}�c�43�#�M����Y+L�t��R�m�����uٿ�e���~{F�d��`�%���3�x~*Le��W��������5�C$�������w��1;���=9 �<��O�����2�Fk��k�~@=qI�
O�ψ\���s�b���r��_C��^9�i�D����|ٖ�M�}���{ŷ�)G�Y�Ac��z�f���^<A�`��+���%]�z�.��i3����V�4����k@�Z�	r�)S;���Vc�y������[h�e�y�`a-�/�~��.	�^�EO��?{k��R�����CZ���+��[��lC#�ۋ�LщH�*a��w�\��xm�E��b�m�^���#5Pg3rpX�=P~���5䱧4��D�|ν��/�؞M¿h�ޗ����p-1��������y�+̛Ȩ����u%�O"���n�hпw�郃=�&6�d��KD���=�>w����m{?}��XW������5�n��x�bL�rs:�v{&m5/��Z�8����B�
֭�44g&L�.c�L�]��ѐT����f��#!e��3T���WU���>dS2W����2swB�U�H�v���uM-32�G��!bo��},H�*(��rYD���^(X��; )���sҏ���yq6+��i�c�h������hTu���Ȯ~�#2F�D�L���G�����7߽�\*��(�0�N��m3�L��U4jo �o�������Y���̨6%N�A�65���6�~&��OG�T�؅����x�p�Q����0T���B���A��q�e~��=1�OOOoZAX�ą�Mr�2�s���4'Ϛ���Z�����a�QA�C*%��k< ��C�?r�Z���GPVGF��l�x��::� 	���]��֨6 Ȝ�o"!�7�(��,��m�ʄ������5�բ.�?��=Z����|�DKJ��`�Z`������ U��R�p�,�����M|�F���$-����Ui�N�~C>���r�<�$�A�?�q����H�}a�T϶��,f��gm��Vt��Ĝ�Nc�;���Κ���j��:mS�ܷ
6Y���I�����?����r���Jr��B�iFJ�\s�];��:��IZ�k����W��p�Zq�Y��P!���~�����$������=�[��'֩vޞ����*��I*���E�����p�TmÄ|� g
����z��wm@�Ж(*=��Jb�D�>7>@������>�םE�g�]��<^�z&�HsfSYs�6q)�R��LID� 4�)`=2ձU�[��h�j'ifTV�	��R[�]b���
	�A'*�0o��(vf���f6I�ov�������Q��2���e������IVj����cK=�9�^�ЄI��jc�l����/� �q?���%`�� xe��EL ��Ci�g-D1���,�/W}ڈU��%���_N�?by�L���b����QJT���V�;-�,�$٦>w�[8׵5o����=���@��5��61���Mu��5�{�����|R��H���������q��)��|#�g���yv�&Ʒ��O(	bK�M�g��15B5�L��d����~3��>��a�>c�zi���<��ml~/�ce�<K���W�8ڒ��ݞn�X~Y?ؙ:`���rOK�()y`ƅ}7�lJE��� ?$���`H'f�la��2P/��mH6����춢���3��5�[*���b�WF,?�V1��]��>���-�#����a9�?=��պ�w'��W$�F���RoU����f��d��+6��)�=�(���!F�������'�m������zBM��Oq��v��-�Ĉ3�������l�Iy!�K��?��?^UZ����j7�(��n�5��J=�ݮ�*��dn�����&�ƓDo�a�f�rޝ�����6�i�1�$�R����l:̋O��W�f�&W��XŻH������~�|�C�1	�1��Zn1���[V+��.ܞ���p�3��i�a$8ߙU�pn}��-�ϴv�QQ��,�$"�^q��P렞��n��?N���Oy#�.O��]BV���T�ۨ��0�K�!��c����Kh�	���p��F�X��wU��p\�8��;�oG}kź%;y���8м��R&�o�Т+�f�\�9لR7�v��Ýэ_o��D:����[��]��(l���yӓCĈA^��mgȋ7Ԉt>[i���S��l�a��`�G��U��khV�0No�\�=,2b9�G-`������� D��u�G��-��]��HcL� R��'��wq�<U����7uŸ�<=�bI��[�.AK�q��E�ހ�� �6n��(�d�Ze]���߫��m�w���}�v�)?�ЏS��l��T�@� �
2o���?4+m�:4cB�9@�!�y��C�1�E�*�8B��Y�ƇL,�5�"�r���}~xWr��E��e�
^?Nƌx��]m��p�
��~���T��V��1���;��a[M:[��O��)�O���:X��kڬ�qP
�
�	������%m�pG�CX��������}��l���>��y�[=L��i[�-��p�nna)#�,˄�-�c�
1M�d�n�L��z����^T�B�RaS{��qEC���R����JtS�?�z�Y)+OHT)a�b$|�����-�/���"���B��#�>�%(��/��g~���&�D��#�L)���x_$R(Ln�b��3yʶEG�*s��yMv���&U7/D��sR��9x}hV�y	a!/koOcK�O��W}�2�?b���^q�� )%Zf@�Wc���(x6/������V�SşTk�7�21������-O����@����4�S쵯�
�w��&���x a!>�dE��'�lP���;G�imU���[<���W����qcZ7\s�J�ؘX�����X��b���XR����Kl8��
N��iA���ď���nɠ�:�+BMW1�-}�4��Z{��/֬-���8h�����,a6>?��O����e�`wOl��
�L[�HU(����K/����hI�'=@��/��^.��mc-V�r�ٮ�\
c�l?��	 �[$"�A�vA�\��y�Z,۟ԉv��X�� v�c"�,�5�f�Cz�TR�,?6Ʈ��zw��68w�Zr��6�� ����Ռ�Zal��
[,�(��7�l���Y�ꇶ�u[���f�7�m�,���n�n��7-�nJ��I�f"�Ӄ�sdOzZ&��PE�5����|�$'��.��G,�4�H�%ؖ�H�r�ɸY�TV����J`C&��;���Hh�w���Ąͫu:ܭ�����#��e���ӵm�](N���|c8$�&�5��!�;�ħ������`Yt:��7�s�TIT�C����C��wE�B�#�_t��Z�u�Q����q����p��ʙ�6����@w)������'�	k��w��UA	�׾�y�D#82��k���E��ZF N�#�3J���Ob�fOD�gc�����nX���@�h
>b�,�C�BK�!�_@�ڼ���ܨ��;��Br��j�U@��|�Ѧ��2���Ï@B�Z�r'��px�}��3����:�D0�41�i�&�=6`WU�^�!/N3������=L�N@]E{�S~w��=G��1g��r|�;�Y��ʜ�>���S�~����>�e�9� ��:ɞ�Q���Y�NN[t�(R��F~I�Pة	�u��&��m�C��f�6���ͪ��hY�~�@Nڱ�Iy��?3��v��@n���v����C����ie5��3�#��O]�}}�B���r����n
1��!�t���h�`Qˁn���_�4�����ᐷTt�Z�>V�:{ڦ��ES	��;Ho&�w���]b�8�
m:�U��؍���x|��o>u��fޯ�g�w��DtSc%�[/�nG�������z���GLr���e9)��sc���Y���d j]{^�^d�g\;���p�ad����B؆[b�{�l�v�ݬñ���Lǡ�~ӫ̒��[���<��&�O�|R>^�<,{��D9"_{������u�S��p�$b9 ��ƥ���F�Bd�*;v�'�i�f5��MJ]��Ȟ������zo_+��:a��,�,w�@���Nh��Q	<?G��S����a�w��v�����������B5����'yF�U�t���+�-ӭ7/� �n1�7�^���;��/$E<��dV��W:�,;�z^e��`����)[��a���d�����S��e ��7и�H4a�|��#�sn��cV�A��ϫ�|*1����m�^��8���$ҾR����Z�6�+��K	��,_���|�(���d�o��p$�h�g_#*!�o����$tn<p�ޔ���V��jPC����hS� %\u0L�c�[�Ъon:ͮ|�bz Le��RH0��r��B�_�������Fi�u��o�~�q8D,.��w�K䳠C��Xq�ـt����իqW��7S��۴��x��.��_��)ȹj�	��ҘܷV��4���1���n�}x�zR`����� ��W���/b���RI�t��L"r~����b���w��`]����S���(�t$�M#���:��<��4r�F�PaOԩr��	Ⱦ�&����q��H��a�r,Q�5��Ty��X.D���V2�][�ʅ���j�Ȑz�+�_o*e�b�m6|��u�]��I­ �#���h���)�(a�������~�u6�>�wgYP��S#�]��I}�K7���0�!JruŊ(ݟ�Ҍ"D_C�E ���9$��j@g����[�\ujo�}o�)-6섓�k���+#���2�Q��
�ߑ���݋W<�w��i�nlܸO� �A_���I�g �	#�ߟ���F����)�l��B��h�bE9�ނt�X0���<��ze��=����qLt頎KH��0�D"���
�nXG�O���nǛ�����u��C2�PJ��
74L��MG�3����͸�~�D���~е��� ���|ڰ�ɞ��x��L��,����P7��܍H�����	l�&#�\T�W)�Ŭ�	YP�_�
X�f���խOaٺ�U@x!�t�VDjKb��.�\pO�W8e��!���qD<�6��>�bc���$-` ��-%����0��ဇ!��b����.E%�Y\ryU/�K h�����
b���� �����l���[!��Ϡ]kp���j�\������ ��9�@"�ז��3[��۪�ku��ZL�C}3bP���q��R�G��V��e���֍��Ao윁����ښ�MF�ai��B�65�p|u���I}^G�B��gM`�'���g����7��&���"j���Jk�X#h _R7ꝅ����1���+��s1�o���@���d�V��+a9l�kK؄�o�&�.�� �PO��
�K$�L�[��-u�q��^}4�I�eĶ,����HM�}�)�o���_���Ⱦ�����<��>�b*�0��83es&�/],�����؊��8{xh�D�CA�۸/>nw���d�@�4�ݯ6e��L��_����cB�XXx$��M񬍞+��.U��e �l�h�V'�m�_�kG�Ʀ���%ۻ�8U�J-ǽh&tW�B���w�I��k@�U�:4Q���%C�yM�s�2&�@� ��Zlܰ������W�U w��Yr߮�+&� u���ӝ��`�|r�R�
�XI:5�x��v��Z�=��{'3I>(�'�O���+�C��d	��)3�٨�CZܸ�L���)�g�i�'��ƙf�ۻ;x�X�
Eί�����r��IdAR��0/|�%�׉B�Eu��f��#%i�@���G��~ܺ1`�~H#?9xXe`~��凞���a��~����Ҝ�;k���)9��D�r=�c9��CpG����Lox^���FOw���̟�j2�aLa�b<���C:�P� e�?��D}�cM�(�t�����(�����SX�Eu��gw�Pv��76���5F��a� �:=E��kQN�Š��l_��ܙ8Tg!���	A����[�'~�[��T���A���!�Q�O�7�@SB� f�Dkߨ��o�jp=Xo4ɡ�F~�p)P�����M�YրSz��0�+`�}�9�
mUͻc4)�Cֈ�I�!�`�T��f
��$�Lox=@[4ۋ���z�r�w!9�`��f��a�d�⊘Z��G���&#dB��1�Z�D��W!�'c���g��C��Ӗ���2�ή�A�,��(��9ek#�9Dy��eJ�j�<Vb�����H��5�Y1#�ZJ/��0�U��ڟ�Ֆ��~��s#����G/k��p���� ']ϣr#
!H���:��_Νg8W�NTU�R�+B�,�:�ܤ���OR~KE+oB�$��R�ކ�bt�m5	�!n0@:��<�K�c�ݳ�G�Tc����=��1�0	�Z3X$�Fw��x��4����q�ZI���_P=�F:���2r%MM�8b�`���%����Κ�pW7d�V�-��jq�	� ��I��+&5�l�q��0�����?�A��!�O�Z�����G�~�q���M"i*�
PH�� ��K�����#k⍺^}|�TD� *A�������O�uF�K��X:��iL�q~�Ml�~���x��r�`���;&
����4>x(���B�U�[�y����kvx����/�ص����ќ�T<����mG���
�^&�S`_�[�u��;�1�:ª�B��ǈ~��a��遏#����̽�.���(�,	�V#X��q_^R��Ft�e���C|����H�MM�"���O�{x�SG4ҦfBD��j��6����מ,U��5�#g�������[slJГ\&5 jHj@������j�X�
N��p<:;��*�$�1� �Tn�[�6����(�}LP㷙��9��)-�2�{~�����F&��%�ў�F��>ªpB�>�Gr���`Aq{d}V�f5�UӺJo>B@��[cI{F&�
�]XG+`M���^��;���)���A^w:QX�-��o�]�!�ƚ�8�%T��G�b��e�����r]��^n��<�鰝�`^l����>�F����5���pC�XO>vQM���Y>�L�)�j?9��Ec"g8������˖���'	Gb�� m5���G�5-��PG1F���>D���jd�iJ����N ��֧����A醴�c���*�����,>ҏ♫����Ib��C-Lo�2�"V����]�lش�+7z��ܐ[8�'8뱸�)ـ�b�5���}��}=_����+����hQ�S��7�;�>�g%��7����|w�?=�vi1~���k�n<��h�F�3�1�{�|�9��ɜ >E�\E���Xbh^�d�x`V�MI������-Z���mC���>˶o�W�纂�u�M5��I#�A�>���8��k���XH�xM	qD����FT�y�4���R#��o�,Z��?˝��3��хs���=&�����O�j��	T�<��4/x\Оk�;�����0d�6=�r��K�Ei����Q��ic7y]����u���: ��ѽ�-'��T\�1_�~Ћo��/S0��I�[5tJ7�d¨��91-��$�kBuН/|l���h��,�P=�����h�!�c�_�*�zq	�+�1(aW���Em+� N�f�%r��ŎQ��"�ُ�W�o�$�
[��W+W���4=��@8��7����5���Q4�ْ���k*'yH��Z�U�)�<����-���n��O�8~���ΗH��3��Ұ��2�Cj62ښ��k'��T2��y�\w��.����bO&&^�'u�	��:_��A���F/�^~�Y���`��,<#���o��1�l ��R��լ
�ܿ|rXKXt&rp�X{f3V�V�Q�=s�^�0�]�� �unYT[�r]��BAgO���򓆓��lx:�^\=�c+��;��lڧۺ"h�(�}�IB�\�&�T��0HK' g;�R��:/�IVu*٫O78F��M�4�}����z��QR�m�ǿE�k�ptX7a+��xV4�4mÂ;���2�c]g䝙�CSf�63�����P���!�Ԧ������	��zo��nX��@��`���_,�G�8[=��֍Yf���Y0P�U����v`^uP��ә�T��lS��#�^�Se垟�%�ҋq�@t��.,���'�
��[��^�<9(!J.(��#/s���r�f�O}Iv��{D�,�$m�Z0+��%҉~ԑD�0u�Y����W7)��^�O������Q���6?XW'��4D.G�vsq"���}s
��{�[���
f\��L��$OPN�W�q�*49�R0XbL$�6@� VXV�m���˸�o��0���8�F���q��D�pC�D�� �DX�G�
�Fe���Hd.nc �H�팇�Wx��ѱ��+����
�ɝ��o��(��`4=�Q����9�T�Λyusq�hv��kVb��U�.u36�)��^�� +.
l4�����[�U\�Ȑ�\M��at�z۞1kP?�=٩���Q�ګAu��ցjY�~+P���J�A@`i�11(�e�b�q&�E����j]+�� ;���.#�󬔓/c���"�VMp�6�ٰ�q7�x<
��_1tІ!�E �Zf�|���,5��H��{���<ѣ��"�C��5�52��X��!R%���֡��2�"�cσ[a\���Q;��0�. �"rӔYS�\K�~�d�Ə��5E[��DBEr�~[�$ɢ��fA"_�R�P��bc#GC���>�2���<tz��#��6����Q����!G.Eڢ�tr�}V��
��s1׸ә�:��@Aͺ�� ���rҘܧ�W�H����Zy{���l@��=�a�Q��6�O=��]��}ր[1cHB(v���t(\B��F[`L�ؙ�<�a{����G�zBiv��o)ө$�O�kY5x��`����逬
 |��i��5f��0��a���SM���v��)M��M�Ig����1��3u׏K��4������^��Q�	p z�ק�uo�Qzۀ����7b�d����>�ށ�� ?dC�K`4��z�NB����e��l�*���������>-��\��E�Ud���&
�o��
4�wG���N8 R��^���h_^>�ۅ��ԅj�u��~{?K�<cg�ҝ������RXio��!U�����La�O�:�	�A��^����{tx�C�n H��m�^[n�bP��~����B�8�\c@�zPJ9��$jGݘ�^���$�qݖM�5�yM�F���L�8e۫�� �����}���pW�[}�C���z����l�3�(7J��z��+*��/-
���%���ܸw����nVp�Am��7I+!6j�f�M��p*�C�>{@�0D���#��׮���a�,P�}+ �t��A4�~�I��l8�m[��H�t�ͱ4O��F?�֏_��9쁵�3���Q)�aWA"
y�\���>L� �g�j�D�SvyK�V���� ˻o�/��Xf��G���0�9�wA�Y��.��X�o������77�V	�(|��
$���=�^VϪ슉N6,�ǧL9)Qnu�7O�f��az��ӕ|IKI~���o����h*��s����e�;�9uU���#�cC�B6bT�l��9���xh�����־��>��>y4pXBc[���T�vΈ˔���6*�����О���!|�����>�$b�a�\}�0�V����0Բ$�����N��J��Z�9:{Ol�n4�L�BB��Q�bn~��l�t0Km�s�ǛT�_C��i��|#�Xtn^f��i=�P��p��6k	�������� ��w����bkN�!җ ��4C~U��`�?t)#0�ʬd%���Z�N�10�<�yC~�zi����S�nٸ�0ޣ:LQ��ğ�b���0a��_�M�6�N���tz�FoL��w�
�ek�~�����? ��w���Ԓ�ك���C<Yy`���A�H(Oh���g��8oa��S��$я�g��/?v�iU/��C�A�C�Lg�8ALS����A"�-,؎�S��~�~��]`�V�=7B�޾�j�!8�ԧd;=S��x't!˔��H�X��L�_6��{C���
�k��a`?��h��릭�U]��Yc�.�9BY� �]D�����FG���q/:/N��QKw>�?�y'��C��	�41���H<'�1\b6�y#	��:3�A�/ >]��/i�Tߏ5nԮ�tU���5��Q���&p]�۪���~����ɣ��'b҅�m�4��ڛ�h��� ���v@���k�N�M߾�`����¡��^��f�g�zr+�Q@A�ƥ�Og��x�+��6^��FY�����2�{��������M�6�]8�7���׹������ɔ�ߓ�@U�?g���\�#�JO���F��٘C�;m�l(�vD>�C��Fܶ��_���	T�"�$��?�8����Q"i�EM���Q$�]�c��+��$��d�4�A)�s_�1�vL��g���9�ޑ��j�b��.��|�xgr<��t*Ox�.�����ۙ�^�t+�b��a�\��A�9]w�)���^�J�u�>�\��z�װ����c���{n\}�Z���D {���7}w)\ >�?�+�[����Ǽc��8�W�ֿ�~u����E�K����|���4�Id��=�`Őw�)H�_I���f��v�#��x�b���L�͌�̾�缃{"�Ħ1�k���q/�	����������5��(�E�
#��H���m����clr�B2�$�HW�f(�=����' ���B1�ӬC�I�£�C���1�h>��5iuz���3Pp� �j�P�+�'s�	�q���9!q��G�U��iC��5##�E�}%�Xՙ�!�Y�P�b���Ru,��	)<J��F��?I辚Ztyy�
X�+������Ձ�hK�_ i�0�f�qF�hV�-�okj[B�<�:��Q�@��u�OC���$�D _����8�mZ���D��aώ��|f�>~)�g~�HcA�7���U�j���e�w�~� N�,��@J��PwB_�C��g���g�s��ku�} 5R�O��ʾ���\�o�⳩��z�	X�����!.� oq����þ�Uߛe=_^v�Ɗ�`�������	_�^R#����%R����-�vU:2jC�A�M��CA���CB!.xvD�|��ȻGw	\zZ@| �:�s1Q�$�muZwF|��,q
�:G��$�u�L�8�xPg���w�DG�{^�X�H'��NUj<d��J\.Ӎ�{i�JȾ���>���Q�JwI����E>:B����S�H��3V$�i�>Aˇ�''��ī��3��#���&w�o%�Tmj�묲eQ�0It����!�O/^�<;�Zë�Dc=J����7�m�C���f5p�R���P�?�?*X��K�7������C��R�y�G a��
cB��;��Χ�b�@��ȏn������O��]0��_�.���f����[N���� ���'�W%B��Q(�?e�rjNG�:�\�-�[�珚���}���>a.]�Ua�B_�T5/���l�S�����ԗ��.#Ҵ&ҒR�+�inw�+��h�R9�p�(zʺo߻#d�^�1`Â�����j~��_�na�0{�/�i��/��(G��-��ld%CNr*Cc����\��>�f��gM�����u!��8��'�O�%��(D0U$1���=�mlҴ�w۝u+�#.,g�ރң]z<�3����f�x롾�m�8e��%�W��R� z�qD����I���x���m��ᴢN�wH� ��W 3[<�%-�GP3E8�a׳X�߉����o�l&Q ��1��ç�y#��dI���[���{쐑QW��P���okr�Ѷ`!v��T�̳������ҋ2���u���c`�Ѧ9���<��p��Y�7}U�͸w�'�m�Ԩ��q�ٹ��dcu�,J�Շ�[@�4����=i�E����]�iAA�
�Xk��pr�Ga��,hC��8k5��LE<*0"P����߄�T��x����o����7�?�w���t�r��/X�90�*�^�Q�Η�~�E�ńm�w�p�Xo��k�,�.�6��'+[Đ�����/z��p���o�1�X��2��<
�����Gl&JF ���L��Խ�t�ۥ�ٙ�Z0�#���H0֕�R�aΩy��"�}��3���2��U�}L���lR�/u>G6B�rRZ��G�f�Ԗ}~��
�q�dF���	]L*���9�ʏ~Z�aZ+zU>��x]H��K.n�8��\�|ڻ:��.J�ʷ&�O�Z���k��c��9��@W�-Bm>����d�1�hy	yzWmY�v�6ck�~#P\� �j~��%bf��~���7�|�f���� � �0��혥7�\\pn�<h@�*j�kF$�l5?�8de̻�M�+I�|Ѣ,�$��~m��K����mZ{�x�~=N�ҋɔ @q��DY�U��e�/北���s%*Ǿ�QzN�)f�41O���6���?�{����Ou���Sk[��x��<���M�k}R?9R�p�P��g����g��e@U��$�Z��i�����L�
������Ҹ�V(zf��%��jPZ*�zD��H�&�s�&	X��AI�
x���=z�H�S��&[���1�Q�I��옡l��O��*�w�`��^ZJֈ�����*���������D���<D�~����n������3F��3|�՗zk+:06��ܽ�ze)8���� ���!eO嚈VQa���N � eq��'Ǹ�-R�K@�Z��9-�9�o��He��QZ�yJX�t򻊯��<I�-���i�G 8z���3�1�ȏ��t����X���)��E�l �=/�_�L���K�����e ��� �[I{)�t���/�W>�#s�G5�TI]j���/0�o��,��r��,�� f�.|Bw��~
X�FBM�F�l;2�����GO���>�F��=����|p�n�J_��N�54�J��wM�q��wFu������Y��R��g@��/x�"[�41��r�/�71�~����gyy���>�F�)�M��dd7���?TAVo_F�����W���'�e�.j)SP[�4���"RD�2�S)C���fU~�imV�wt�M}����5f����ْT�Q��Z|Wtj܉�r;��_�bn���G�;�Py�~!2
d���N��GBkAx- FP?����򳅕�G�w�j�L8� �崑G�&��1z�t�#H� *@O�� YL:���ݴLR�sO��%]�OB�# ���N\�<����`��+���گ�7
؏�C�4�%l���)$�}1�'⯰M&uĬӏ?�x���s/�
����o���,���Yh������������n�N�`�F���/��i{9�����'��_
���P�������� HU%�!�3.A�P �3�b���*o�1�<&Z�1�lmv�E_f9n�2�O3�LG��q�6	XP4H>��$����zǋ��1gN.
2 4����P��	p6���c�)[�I�<=�n��l/2FЧQ6��Z�s�yw>��0W��T쥖�m*w���c���rsmaI~��r�a�N���M�mS�1L<����b{�I8�j����5&S��K3ܐ��?C�/��S��@l�wmR9� ��$j6��3`w��2�>da�x��kN��L�?e�����]���5��j� �#�}qG���M��y������T�%��Hф�V����K�����[�i���@�09��-o��9�����
�dS�GfՓ�K��j֩�lf�i�F~��ހ��>ǃng��OkFM�0�#����� ����Z,C<ɫ�Ԕ�q-씲V�v�} e� �O�*�0�xLwj����Hw��#���"���Â���H�|�oT�~�)"�T����8�ӕ>s]���Q��u�-����w�W�B���is>z�n̽���:nE���#3�vV�cW��>+�7�\%���>?{�>Ẓ�kj]����'���-"!5����sf4DR����7��5��u��.f�'���I��ٖ�)rM�W���)���D��p���;�	�:
����:�bm'l�� ׫�z�퇯�%�����B�?1��K��9��CM� !�����*��S�%po�k`��J��
�<�,�x���L��70�ҵ�sG���5"�G���o�t����Ww�8�#q�Mǌ��/V/u%imo:��3�YC������oC㬶��<�;�����E'	<����-+ܼ�\I�_4|�y~5n����~F���{O�v8o�7� @�P�fB@G -!��:@W0PTd�eC���J�[h�zT�d��! [81�C���e��Ji��#¡+3	9�+�I+�I^լ��o����RL���_��v���C�,�0����ጇ�-TFH�U07��1�x/�A�b�g��)Ѥl����7������2!ts��}�P-�T*��6�V;2��di���%g�V��9�*�.Z���.	�3��:~��Mc�`�w;����7d-~s^<�P<�)}�"�p�1R�W8�����!����Zc��i�m���j�K���&���n�b���� TP4,�әx�ߢX�`r�&4���W�by��y�c[#�]3*B��C����8$��@�/C����e��B�0��x^��f��F���A�䶱�d��ֆZ�!�� k�v��0��6tq��M���!"e2:�X�p�T����LW������X�c�q%��^Y��5l<%(�64q1,�ؿ�%xu퐇_.�&����W=t)G�PX���6���s���k�뱨F����M:~"Z �|~�_q�M�R8�z�!�z�PI�n/��O ��V�d�Ʊ�L	AN��hy���̒��~��	<�����a�Ͽ�7� !��|��$��ЃT��Z�N�r�2�$�z]��Q2qO�X�zOx&�$k����A�$4�]L�-�}a�Z���m&�!{CA�;��t+ĵ@����zq�����(��3dl�c��{�d�xx0?�yf9H��+i�wZ���|/tPc1��5�
x��U���D���|�0� 6k�/Z/^u�}ߖ���p7tmQ̙��?UY����S��\.��]J+��{���:HH���3���||.]:�D�'��NL����;g$�
�#䏌�ou���JS�6���B�,�89�!�)�U�z�r?�O�N�D��1ƀ��<7���Y�����}�*V�.mrGsZl3o��3�\8��;�y�`QM� rP�Aύ�7Bި� �b�<qH��+��H��y��
eq\> ^�+vEΉ�^V�3����/��6�,���z|�����,:NV-�����Y���9��#�T�r�����d���eש�X��KU?O۟�!s����C�L���"�ѕ�R՛ ��r@���S�@m;���k��],f�C{oJ>�'��hl7	�Fƌ ��vv߇��"A�v����d�ѣ��ͦ/-bH���,,1�6+΅��)��^��O�)	v��~e�e���'��n18��AeZH��������p���0�_�
���/ʀ���bhh&�~a0|[��]\X��VHX���0&z��7�NPR½G_�d�șG١�q!;�ۿ4��_��Z@π������=��Q�v���Lћ�>y.��g h�w�Š[�6e1w.
z=.���{�F�F����� ���J㤕��2����C(��v2>ڍ�SLҸ��-����0�Euoo�'�F{}��O�n�p��60�ig@�$�r�Vr��U�-�'���l2Mxhȼ�����f̳�3A.���7<���m�G���_��[M�7?�Z���/8R����䶥G�O��;y�Q
:�Y+*�b��H���t=zt�QRiu౒�TZ��ùe�E$V��U���?��9A\����+�A��Qa����3��PS���Ƈ��Ŏ�B����+oR�@Kni��}\�G��B�J�=�ұn�oC1�\�QR���
v]��ə���~���+h��K�x�����d��0"\�3�Xlf9 ����W�㱆9sܕv�]�p	+H�U�7��2��8���K6��f%��#D�a���ȴ����o�vEec��f�w�=9����%9��q�Ն�
r� $�$\��j�W&�E�U���@t,/����4(���H�E��t��7���)�
�M�m��>���+�<G� <O�N�G�{�ĳ��l�&z"�	�j	��	������e�̖w�M��\ͪ�q��!��}2�+��
���@]G�L�u~)���E#��-�a���AC�����NI�c�����E5sR�c��Ni+�<��n�f��}��I��'e��TD?�:�`I���%�T-.�/w�-~H𙄏#���B�I�O��/���m������,�=��c ^�3s���k���;�}PI�>��>;]�=��ֲ����GP�����
�������i��:(u�+~=wˉΈ���BU����f2�>xt��b�Ln�z��7,4i6 �� ���n��,$>�P,3�3=E�{]R� >����`��<�/��e^�!�Q��_lU2��,į���3X��Cc�<V��]h��&Z��RЀ�u4c��2y}��*Uۯ�EY�%G�=-,��R[��l�J���ʕ�{�|�<K���os>�.��546��ɆY`���?p.���
U��ٷAw�@���E`�#�*�2��˲9;h��'�d�VS3�OW	��<},��b %0C%���걇%�fhZ�YI�:S��ޯ6�i�p�Img�D}�
CQ��	��UG�qGX�_@Y�^Ҝ��r�>��@<�O�tns$tb�%���v%�\� #�wՑ��Y����tӤ�Zp�mW��}�u-I�b�!|�H�X��ʝ*_֞�1a<�fg%PU�Or�ء�L��$�|�P��1�*���"mif\��7ᄝyC��v?�s���$�aJ>�v�KT�=��a:Q�X+t*;Cb�.�~��6�c��/=�I���������[52��/��Qr �0��Q��R5W:e3[�%���g<E���;�k�ً��=\�58���o�6=Q�?��Y�L��!6x�J`Ogթ`��o����z��}��+�/x�O~
K<jX��,�T�W>��|��=�����e#�Ki�nޗdr��D{����a
�m�m������ѐA3�6�A�2�Hm˓���&k�4 2�w'�}&�FκM����ډ�ɍ����5C!x��U��t���AK[�.�]�(=h�H���h�D�5�/�f�Q�Ѧw�9}٨~����ܜP�G!۩�a��{︛�6c��7y�pl8i���ga�'4�RY��mU��Y6_ܽ$�^��2|�9��� @�(����?K2�M�Wʥ����qWw�JW��v��\�~sH;�B�Yܸz��4�HR�rS]��;R��{k(^K�\H�Şc� 
cf���"���2p���*�f'���t�;h�� ,�a�jպ'�A�8�)��(�6~[�x6�V-c"r{:���
�����,W�yɉ�1���g�e-ꚝ+H���=�Z��׎.�L�[3#~7G�Y]��ۓ��I���bFA:#�H&}�4�B��D�)��Z���\��
��߱�,��[���2��ɏ".G,��nc=t�|��z��AY�w�1���e#�̶<|A�6��W���9qA�m��D[^���풭KVק�s0|X{d�w��m�{�c�f]�N��y� �U���~�GG_6.����|��z"7�����\���H7u](�g�4&�!ʤUK(�b�笯�4!��v��P�����������j��SǀA2���+�>z�g�^�U����1l>��ɦ��h�c�+���+k$#6�$�D����>��|`�����!���6
�~��&��'�����fnK��.(
������~gV��G�^��g��DD���Q��Z�a�$Y��l���Qj���� ,�}�d#Gz	��y�AJ����\�z�:��XHpy��M��n2L�˅^�v�wk-����e�ǧ�2�L�����e1�ZѤ����+0�W�J��� 
�W:w[B����3�̢zU(�[��TE-Dtn�s�ͽ��w�nWt`����w�y/o��`�����][�� I�#�����܈�^P�� �,�5�И􇪊�����bt����鳏XS�Mt��2H,C��ή�^u�6��{!�Pw��7�f]��#���ޭ%K_P�HH0T��h�������c�	+����� :�+�_[����a+�l��G zv��s�I��tk����\����/��Ep���)똭��
t&1���n����Y8/���1үď��Jw�TR���M%�T*J"�����	1/� Hݣȅm`�`i�f��Ti���Ðw�Y�C�[���1Y������2p@�O>*DJ�߷�V�."���i�������hfu>@������t�"��@Ů2��/���)�@0�H�	����H�|HJ�]&�0�n��AwW:7{%ۑ���n������_ҳگ|���M�;���ۈ.�rag���w���t��D�Ӛl����E���w7_���k�@E!�t%�([aɂ;���@9>ꋭ��/8=�q.Y��,4��	��غ����#lv����(9E#��^q�+��,V���!J�
��g�ZD��$�%��L\��w�����W��Ã[I�BU2��l�d@;��Dmj�B��n����������@� �mk�N�%�έW
\���N�lr�V <ϓ���j',q��?�+i��p'CF��\�����r����%^7h�+���<t��g9$���c�t:�6*��A#��{��^'$Q���q��x�ٜ�K<;x�����T���<��5K4Mye��6i�̦y�v._�����kK���h0T�f̰w9M4kwmw�1�"�pc����3����`�Bۂ�
,�+ՒI~����l��`�]Qd�c�R�[yM4�6��wX���$Yc�^%�_�M�u
�s����r1��NC6��xU�G��
�m�.��	�贈�V���:(���
j�K���c:KȾD�XT=������m˩��8��AX�#��#1�c��Ehy	sb,C��(�I���v�yO���eDu��P4ƫ�L��'��7!�0p�e:�"TYpV�D���`�F�	�Ȫ�)�Y���о���zFk��}��h��0*��~�D�����31%t8���g����ڴUնش�R�GWA�[���+��w*T�$��oly�[Z�z��y�x��.0A��S���W�6��޷�����U�q�yz������Ԯ-�X�sl��e�G>e�a)��!���(:�5U��6/��H���gقQZ��}�z~m�ZK-+j�z�h������~2�����U��<s���|�M�aHB���!S�!�RFs|�?7	rщ֛y�&^%����֬��%k���X��|3��PKCe�05½-p�S�͇�j�K��D�����UhH�~��U�>=�� ��xO�4�?.��w�E��k��S"�up�_I�u�Cu�Z��$訟h8���x<)"��Y��䤍/�~9(�����`0:�r��k$R2�Ύ^yQS�W�ƀ"�	��.r��BS̬�����YÀO��͡���n�:�
{Ի�[��&��>C���ݲ�Zi�	��bM^8��9p���(��z������~��-�b1z�$y$�t��ʐ\���uظ�x���;�x*
��*�{���M8<d!��mpa hcT{�+�l�]��
����q���{dK�`�7P�Ҁ�lx�el����Y��&���Ni�8��u��fEm6<y�R12ԓ��#bd�c��X*�hҕ�+ǟY	+O/��
����#�q����Θ9ȓ�PWZ�A��ji>@&ي�M��܆&Upy8%���5���{��Mg�����}���p�ӶE����7�⫅��:�6��}ǐ����Jȱ�Z�, �6��:Cm�l�j�����).b��k�I0>�ybw��%�,���DV��}��ڄ�K�7H8���\
�2M���tl����w1b����*5zЃ����\1�0a����ƌ	�ǣ�r�V��*��x��M9��<���v���x�/���8#�UIo`�|��f�W����}�Ͷm�У��<k�������vh楄�i���w ��BR��^1J/lqɁn�I�k�ڛ�M�oU�Ⱥs0C.h�<g��9��R�+P�������f��<D��|v?��pe˹�fv�ݰg0t�*H?��y�J
ϭ��8��2k��&�b����G�r'S���o��I� >LdCq�f�K���@wک):�G@��e�L$M�� Ǡ��?��Vf���x�!E9��vd����~}M+��R;�Ҝ��(��F��iYd����.�mIj�D`������(B\��'�hT��#h��5�?U2��`���=X$��jv6�xp�w�e�׵�r��'���Jh�̳�1A����c�6�����]���$<9�i�ܹ��5z'��ԡ�эE���^�˯	r|tf4YBeG�_gd2P�&~�Z�d�
jl��#��jp!:�[��4�ƒ ���k�YG.Qs��xӍo��ҏVQ�TNl4~�!0��<�6n=��tO#�!���q���h�	ḸOH��3W x��&�mD��4�:cC`�?�~�3Q��6pb��?��ۜ��������
2�9���]�"�;�}�g��G0���b��K�NKD;f�2@
^���p%��<�z.�݋+0P ��;ˈ���x�T9f�o>!��4������D�m!�+��E��?�YX�_��f_�Ȇ$u��(��G

X`Ö�QϽN����?�:��y�'4i��z�+��XV��H}Z�$���r/(�򗁇�}uGyzz�-7c�R��<t:+�[>�pKW~�������]ײS�:XUBhK��.��@t,1o\֑�J.<9�-�T����4���}:�"��['�
G}�9qz?����3����\q�mϸ�g@Tih��j��$���o�w���!V=*����V;oSb�TL]ĺ��JG>�L�����)�HO@����N�&r]�w����&#����,�%�����)Ǥ8؛o6n�n, ���)��B�^�5P���+���:Щ��9������Dbcfn�a)���4.�����҂��UH�6�Zfڥ̴K}�T��������]����J�A)��%s��U��=p�1)��#ڨ:�zx��\��cp̚�D!������Xw��j	E���O����(p��( ���n�6�p�4�G�l �7o/F4w?��L���9ˌ{y�w��~�ЙyN�ه�Epv��'���?�``���ޥɗ�`����\8���R��R�w��&���v�=ﲳ�u��#�iE0*FvI�H��bW��#��9C�,�
���dX���,��y9���<F�dWx8�`˚&��&���,X����*p����8G�G��ص�������Ғhpe/��z����D��FS���G�@�"G�ͅ��܏�����o��)2-����e��F��H�G�� ��xu�[ �:Lax �p�{��7"C.��I��;ق�u׫ mF5+>���a��\ˎ�d���Ɣ+Z�a`�Wb1`.
���+��g��G���2�?�$���ta��ց��"JT~:6G[�"�N�'�����ׂ�����w� S�����sK��n����\�&��>��݆btK#��2�2m���]���,���9�*���jbl�ӳ�u�P����{���N���E?��(�R��������HvA�wa	��cս���=��J�	N��A������jSbQ����ynSu�ҬJ��|���D�&�O$g�u��>�ռ�H���Z/�u��+ؽj�J1<0Ed��Y��������fN%�^��{2_#u�1������KR��(�o��&��3�������u���[���� =���\�e IɜL��"��Ze���}�G8e��PL�u@!�_,h1��l/�X5�M5f�+l}�� �[F���q��4��v�f��:�nl���\Sb�;C��Y�vDQE)��[���4g���y�I���JBW4*��)Sz功����+&����g&�MUTw���>�9�� S�K�m��%STm�jyU(MМ ��q����NV%��2��S�L�Yp;��Hso:�����m+=�P��CE�'8@�@a@t��aNF��Q%#_� �K�r�SD(��
:���b)q�bL�eА�Hu{��[;]F�QE (�7��8�hNV���'e/*L!�q�cYT6tw-�5��_b���yzr3��y�5���Z��,���X͒���e�L��	�	�;��Z��Ȫ��g��HG�>���`Q!��ҠW�qtE$���_�)�0�D*mV��}��'t�ؿ4��y�-Z�d$&eLc}����b�c-����қ���ݢ���w�ȓo��6 ��Wp����. �=� ���ˁ!� �h��8V��D뚙b��\�U!���U�#�i}�b��IHW�Y.;�%�!T3�[ޔ*o�_һh�(19]�uu��|���oSѬ��y�C��EFL�s�|!�=�"�����E��=�~�PHR���`���ˊgi'�ά�S��l�x	<0�=�0f�?*@��~.4I<�ǖ��g���K�P����_��Up�_ƺ�`%��6*}*�j9��S�B��C�����!:1y)<�{���I<mw;��|*c]��VZ®�A`����s�=itO��7�-�Y?z�~�c��mQN��Id��0ػ �D.Wn�j{2��&�kLM�n$Ϛ��S9N��?�`7c��!miy8M�IT)ӆ?���(��s����A�s;�ӺO�b����L��&=�7�dVGs�}3���^���6��(ԕ�k���կ"����\�٭+�GvŔ�^]\/K�N�E�C�_t�����>�����{fC�!�ȆGӱ� ��mg�^�V�|VL9.z����t 7'P��z*'�&5����'���k�v,����U4ޓ�B�j{��c��ߩ(���uɾ�O���$�ItD��>�v�g��O�J.f\!0+�5�!�$���4�h0?�? A�o~D��"���	��Y�0�}��}m>I�qt.�A	�V��i*5&aS.ڿh=�����^��f�v�$���+A��i��[IFJ�b�*+�Ut�	��w��X:]�I+#����k�1J�F�m���ĐPJZ���JXd��<���<�b]�l�kJ�	��-1Z��Z�
�����;M�1܏�ْH�D�|�Vj��JQ���!�1��~���S],)~���K-D�x�����EI$
�<{�o��M?�QZ�XoRV|OVǮ).�r}�&�&��0԰�y�}�':~I�Ć!����q�^�`���%O;,.:&������:6�c(�Q�ޞ�s3K)�N{�E���I�W�ÐЪ�J�fB�R9� ��#�r����ӟ �e�?Y�f*b�Y��*ل)JOYU��p�8�$���:���k��RP�>��|)���'�,BQI�~�I&�:J�7�Hw�K�O��B��(�o�/XP^a��f��
�5/�Pk��#H:�1hA��ɶa��� )V��WŪ��7>|�,*�V+7Ȩ�S&j��H�ڜ��J�S����'5�� ��^��t,Xd��oi�1 Y�9i҃�BU�|��6��	��('M�g̐���6�0�R@6�M��N�@Ҕ���b�G0[��S���gr��cf�;�Ȼ��]"��m7Ȝy���g�}��=��2�?h�A�
�L���:v������(��<��l]d�����e�va�mҟ�v=�^�䉴�>	�e�#��Lv2��^��"H�a~V�����,;��e�ӆ�4eE.��#���.j�L�V���nc"F�/:x$���O�i�y[�9*�>��]P��R��,�����Ț�[^~�BO��-�O����:ې�,tQBW?�Ϗ�g����iojm�晼s��fY?j	�P�5Fc;9%�˱_��+��vB�j.dz~�*u�x��2Q�SoN�e�3��qc|/t��)E��&(m\�hυr�ɝs�����1"�D����.m9|Hn�AAο��!���D�[";ֶ]���?��ż�L�U���&.D �8� �E�K����rO�q���4#�~6ۓ����램nb�Ia	���j��r���:HfK��Բ:0��׉Ƭ�r��c��� +'
�u��Ay�$�u�m����G�
���T)���Pj���!���6���w4{����s_7�0�x3�&��a	��H�����_�ZF�+���t�'04uǆ�����|�
,B�m����iU�/�b�:u�R�r��[�\c9Ûs�s6p1�}֚�I�����v�ĢD�ц��w�CNiY�4�\��q��볖��įDNpA�U��s���y�pq��m��}�U�H~��۱����	����8y�.��(~{0�����w���{ƶ������{[!��C��u��6" �~;jf9�&Z�[V�/ vOR�r��t��a&c*�������=�=�jŝ�M������xw`��a�F�Ҳ�jf"�@m��b��R����<�ՠ
��?T�ۥ�%��S�]�.z���Z��.R���p�}��d!3r�3H����"yόг�bPw�3%޹4��
J`ߩ���sO1�3u��Og^�dE	ff�I�����Հ��k�oW^��*�~���9«�#��n����-�	>�*��l�k�Ml�^�����0z�32���iO�g���s�V&��y��v�=L����я��&����yx'�G_Sw]��<�W��R���E���`��&3����G�U�Q��Fa.�C��(�iQ0�8b*�&���d����[c����/��#)��@K���:�ؘ!>]+��t�q�"~�bp\�%U$��Ob��a�Ǿ&�H�=z����D�v{�]�d���عvi%�����>o�ŴɌl��37$���)F[�t�w���x���u_�«��ذ�VC���1Ĩ�1�~�v�ﴍ�0�*�3��zx_��]}R��o�����t�Ah�Q6�V�����/)���Nv��)	�h�����rD㔍�Q���j4Ĵ�u��g����,�B�Mқ�똳T���;���ѾV/ ;y�:b�]�:'C��	�=��/�䓴����~(G�`,�8�վފ��@�I�<BP�����k�F��Z�{�>r���Qq����!'`�{��
�k3�3��X�$��(�G^j��\�=�*P�*>z~���a̫��z�ۄ��*ןU�,��eqR&���W�d?���[����ƤJ��2�k�����x��N��HPvz���Ӄ�?)��y��R���z�H�CpB�Ы���w��WH�3�ź\Z����6��V��B�Omo��V>6�tO��!=��jZ��ywn>G��<����h ~�6H�^�>V�I�Oh!���
g:��ϝ��\�f������>P;`���QR����I�%�Ӛ5�7�L�V�!���:LJ��yG~�n��5�M7�giv^�s���4U�' 䩞ϕ�(�'ío���gb�C�%��M�j��P�y���`�Q,�>j_U��i�hhw��W�Y���}E��6�%�Iu�瀭E
7��6�v�� ��E��G4mG�v@O����8JQk����B;K+0Ǟ����#��ޏ�eYF�T��B��t8U��]��4��'�t�>V'C}ku$��() �4QD4�>����vb�_.W<t?9.a�8V[c�P
z��Íط�����t�@w$mϾ_�'6޾!�N�B�)�S�0%����.C�)WO,�H��Qi�2mޛ<3���K&��[�H���/��IgnM$Jд�6^��CZ9�a�l8������񝧟mf��u�hr�t�'�Gx�Q��J���>����3.8�}��*��q���6���P�R�y����ڬS	� ��ࢼ#dc?�o>X�"y4�zA�,�j����j�Ƌ%��nG�>U�t�k�h�dYT��J���
��5�U1ֳ�>V���iT�MO�^ܜi��Dĝ�l�y B�u�� �T	��|Ѫ�d=� P�7Ut:�}��<�?	<�������O�Wut[kU�ˁ��v<<��ޡu�9F{'�yWb�:���)Q\2�A��eL���.ӻ]♴���kf��v2N"$�	��k �Rz�@������TGhWg�j���t�����3�?�Ph�t�	��2�+ɁⓊي��=�]`���s��	���[��	�ϑ��2#�6�}w��M�6ԚdA�e�O:�ފ��̨���M}߬]
�>�0:�����պ+���i�����27G>px��HO1 �����CxM����n��Z�g��x�$�X�[zm��^�,�Cֳ&0I��'�Q�P�i������H�VU�vx��Y䠏���|��/x���н݁���(\TH|���̪��^-�vN�C\n��*��d�U���2b"Q��3�āB�Sb�=ç��s�����gDNC��}�Kl0��X���,o`m�<�}��VwM�?�u��'4�ݕ������DoY��RR�pQ��3N����oV}���K�}�R)�c�ǻC��G �q�'�}��J��7��UD���~Sj0�LcA%) X��~���=T���E['�ɫ*qD4����8�ŋR�A\0�N	)�?�e}��\�����V��*�1@�_�>$y����z�匿4[}`��h�nv�D'��B܅�;n�Ia�݀��-��A�u�'`�$�������
ާf����#����R��Bs�Iج'�,�A�c�=@�'+1��*�+���2����̔V�,6'�wEU)$scx��D�"�:� �+��
�Ȝ��K=�5�mK���ڠѶLd�,�i�V�̙�iQ�Fϝ����f�v��I��T2��~u��=���wJ�s���R��`��S���S��i#��\��âx\���jyʊ_�xye��z`)�̰����Y�Hl��R=~T�{����;�!��3��7�/����)\8��%�����ʷ�)���h���P�G��գ�E3A��s%��M96K�x�h�}���`���0�sÚ�-oƈ�'٠w����IzZ��La,8��V����)�H���=:%��+� t����`ᗄk�)���R�D�d��T�"����ڄ51m�l�)��Gs�=I*!<��T���~���B�f����J
��a�h	;
AKǙ�3B8�0��B܌`�J%��w���lգP ���X�7�����~6&[#�w)ύ���9�i2wA$u�H*�?�bTD�+���Nj�>�28&��Y���fEpsv	qtk�閇%��B3�Cd����K%y"`�"Pp��ޡ�ͨ�M�Y�o�Z��vGE
��)����V�s37ϫA� `l��>���x����Z,�V9�X"%�۩M\L8�v���Š���R@{�Ѣ9$��	�1��|;Qx8�9SP6E4��xu��[ߓ�W��^��t�v��j����t�GH%%�މ�!%.��w�`��N	[�h��@*3����5l��s��M<�WL�l:�&�:N��NBob�1gq&f���dr�f%\�����Hۈ�$�Ǟ}]��"z��.���NBQ���D�X�����`�ߘp(�b[�#�Ja�!�;��"9[��I�l�r��Q�1KFUA���qE�³��KrtA@��<��lz01�	&��p��lG@�3cG�x�������E�����М[��r�x9\,�5��S��h�J��u���\��������_�w_p9�Y��9]ݠ�<*yz�b���~!/ۢ��n*qC^��#S�[�<��r׻����X���5W#-O����L���.��
7�pJ�0䉩I(L?����I��/@^6� �ڎ�������r�5�UUd�@	��Q��u�㸛�8ӡe9���t�"n�9�J�G��~+�Ч��O8��jm;<�4ъ��bI��w�N�)�97G�P�n>;T�ᒖ-����4����9��%I4�`u���`�v;a�ٽ5� \��(���N*�M�J�r��:�M>a���K�A�"A������y^��'�B�*�lGG<�R�Q�1�os�v�j��%�x�\��	C(����<j�x��+��uz#g���x��j7@����h���t��}Q���]-B?_�/{Y�C���v�Ȧ%�7Ϲ:��h��	ϡA6�p[BUrٍ�hEe�nM2��6�-A����e�`.0�<q�
	���g|���8U�&�gbW�67Ӯ�^���_����7�����;��5hY�~��}�!8l�*��y6��Ke�����UY���(ʜW7t�T���*��.��}'�)�R,�b6���r�z�0 ��B�/T������[��>ǐ�t���629 y;���y�e��y"�w,�{��3�M闐p �A�5�Xƣ�o���ϱ��<��~��$úF��
���]����	^'&X�������'�LO��R�ٷ"��]��Ys�d�WU����v&��,g�
�aS�2X� �7�B5A"�y�\�3��I �R|�2����sx�,8����Ld��c��i�1X��	�4�z�yN��p���έ(ǎP����}ۢ����)�'�Uc�z��?_�\-������_PH��4(a��;�����=*��Щ��l��w��V�*����yb�"H~8�Y~ �� D���k�]�Eq�%�n���*e9ZH� 훈9Y��a_�$$R��(�	I ywe|*-�_�X*%�)�0w������
�l�*���C�|fo���̫�=��J�����Z�k�缣��"��E�V��./DW��
8�K\�E2�"-X�$�L���2Gx�@Fno��04�>�9N$��hA�V�| 9B��{}Ն��3�~�
��6J���t7%$�=�pܢ<����.��iJL�E��!�����	��X2��8 ˚�%+� �KՆ$Ϧ����ō����M����d��
��T���.�ؚ~��}�)��#�H��P�9�s��ykT�����N�"�J.����N4����S��������I�C>a��*�ӕ���}�ok2c	���^}a�}�^&<�%Z���D���w[�[
l���B]�� ���oA�F�>k�>K8+����\�c L�( �� 5��`�pk�Egf�գҐ���r�MK�{H�Ӎ�W���Lf�y%�+�c�w]7����n\�7�$a ��x/$ɔwH����G�\�A����鷋|/���↨�x�~�Żk�O�e}'����\Z�����a5a�+�m�[����ä'����ZVLC����95E�.0A�m'sr�Im��3�]#����/KՋ�3~��Z����Y�����C��A�u#�⁙���i�0��[�`�Ɉ��"*ur���Km�������e�3���,��~���@ �P(�%D~��Vƣ[�t/Y��ǐ||���ܰ�y-Wi@$�`�V�j�Z�����@�h�k�0�u�lr�����+BRq/�[٫�S@O��33�v{:�Ʋ������vAWU�ǫ
]q_�#�i��
dX%uJ����z!Y�"� zmȲ<a1�X�`@K4�`�1W����1��[�R��!��@>4��浒�,Q�6�O�>-hCI)��W��5R��@� ��z�PiGͶrH/�M�ÖJ:�z�\���{�#7� �-���w�s����U��g�i`�������v�:W�{cEL����q�j4Zԫ��z��U�ZQ���)Y�7h#��u�)��ߒafxe�B���'Ҁ�Ý��-M`�%=p�㣼���븍��#�7�F�L�����N���ϚC��<aY���e^�S+�g����a��c�B�������t�l׋z������!�Q	�ݕ�+R��r%�k(�����8Yluk�E�0'�b	P\|�KK���#���{d��s�_8����c��cE��D�!�[�����J�d�\0+ߢY�x���O�[F�#�z �:f�S������Tg���2 ���I�
�U�C&���X��D�y§iBO�O�54�Af�Pљ)<٫~8�<�|��I~ʲ)�Y�ҟ��6�@��j���T&m=~yVƖo<�x���r,�O�]B���W�k(�)�35"42�oc�8�+����N?�������j�5
��0��h]UuKģ׽�ޕ�[~�#�-�Δ"���W#Kd�/� 5�|���g<�����8*�Ǹ8��$4����d���������}i�I|`�f$f/3��[��\&������/������qtp~(!���Ts� �:��ٍ9�6hy��Q��$TKuP�<h�������=��@��kv�=7F� :�6|�ƃT�-e���p�v�ڿ�0� ؘ�9(cg�:��Z"��-���]\=l��FM����Յ	�s&��P�pQwf�Z�c��]�]�p,-atј�Ϻ��	���5��9���5��gO3]�� �\I^��-	^c�2��@�[q�ɰٱ��a�z�!:���ƨq}�� 7���Pr�e�;=�A���=8��R�����4�o���(xcA�\�=�)�NW�B���p���[���\�<E-L�2��#�7�~8C��X���b?��.A!����.1].� ^�b�}�@�N=������/D9M&�V/��:�0�~ %wđ\%Ӄ���T+�[�Q�Z����"�
{�̺f��t������F��ڕN���w���N��мgz�k#�a7���87׵^DґW�'L��]
��4�q4����3�|��m爄Q1nˤ�
ɐo��%W9�&��kY�)�5��}�x`�% lm���ɪ}�Y3�Gi��@蕱%��n�)Wb�f^���b����C���rO��aV�-c�������.�h�m�,��0��NĒ�K��T�4n��Ҙ�X
!�Y��˩�r`V�$d%��=�NT�9�B�eT,m�)P�˖�S�(����"4v��N��w�'c��g!�.'�ILyL!�Ƿtv�h���a'�;�r��.<���ѷ�hu�"_����T�`���p�-��/�Ǯ̤��
�� |�S���
c��� 9H�77��.E������3��? aj��鱔�~��`�˰��m�� u?��.�=��6}H��md�{'�%����{����R%��IF��&�*%�(���oPꦽ�C�������QEUՒxb�Jyg|����ef��j M.˯:\M��A܈	:Sp��]��H��[����&�����+rV*�R(�J���Q���������?i���I���kJ�v��dM%��4�h%�*H��y5����'ʁ�i���Aҵ=��I�7��p9Q�V�o�l�6���4^��CvP��x2�����fߏ\�(��L���⺺	�C�KY���h--���I͵��Qk2z;�}����s/_e�zƱd R�cJ����n�*n*�){N������(���7t�V{�c#=�O�L� 
RUY����D�DHa" QѠ=�:S0�i���/�i0��dj�h"����N�[[��]i�����i�cx<\�fhB�P��UF�I��kE{?V�Q7z�㈟%\��
��!g�s��ۡ�o�A�	�s�\�5�d�hs}k��Ԧ���,_QRB�` ���W�t�#���9}��A���ӳq���a��9P�a	���Er�!�,V���H���O9��Zz�Ќ��>S�2��KA��rB���d�-�v�J��U��y+��̅�X�r�Xz�k�}��-Ɯ��_mU��LT-K���E(vi'g�sV��;�f�@�+|��h�`Lݡ�*�N���Bl�m��Vm�n�;���¼
�bf�p��)��ݸ�V[�5Ě{.��Ě���т>���.�+Ҏ��G�E)4�x��:�U&��4�*���v�q���|$A�Q4r&�>بo�d�rP�R��R��T:w���[��f����=�zo��h����O�[Yc�{/)��	ne��RE�͉���ԟ��q�(ٙ]���Z��C�9�kM5VԇB2���{� M"ub"����-����'s<	��,�J�c�j���1k*,��tL��u��]M.��Lb�5례�^9;�"��ׇ��څ��� �՚�Ӊ�\�=��F�aj�޷��ˮ�j�Ș��}$} wTJvZ�XtDV�#
Y�e]��K�<���o�.��I�W]��t;< -�WL���j�G�S<�Le�u�Lȇ�k��	K|�i��T���V)F^{�=��
fyO�W���|�D��o蹹���ԕ����?�1���1,�)���@������gv�ɱ룓
���vj��a~�n�.9��&�ݽ4�OJ�p�V��f3Ʊ:.���_'H��m�O��#"7ԋj(�l�K�=����{!)x+i�~��CrSօ��X��`d5�Wm�dT�z
���c�塸��J��.
�Zܰ�Q={2|�xtn�����x)��mT�،G8}�~�K<���u�����9��
�o�)Wԇ�����8�<�|���So�\�F��3tNb��=Z�=��9�3Z�E���T=��5��I;ַJ��Fn��p�(i��p�E
 �(io�^?<���s�C̝ʊ!�`��zn�Z�U` �A���wY��NA�'BEx1��{8:QQ����m%�f�&K���+f���qwʅ'ҟK����o���gQ��H�ٗ'�Kʸ=�BzHM[P����n��� �?��\��-��W����A{��xm�<GʧF�jq�@���ް�t�Z^-P��d���wL��>�U~k�:�'!�Ň������d4F��|^n���ð5=��\	�ޅ�*�������!� 
�����um��X��g~6pQ)| �B�'�[�F����n�2 �߹5K!��L�E�셷�V�h��&�L9�=|b���rJ,%�(Å򳿑�۱�Q4���l�j��$&d�.��'��t��ѥ��Tڬ��?��l?��3�f�3!�fM�1���*��7��#����X�L��Γ #;� ��ڞ�7<����L]���� X���'���TB�&��)H�@;�ޤ���Hʹʟc������#gS�*�� u���5��L,�^,!�W�� ��|jM�u��C�����)������1 �p�K>�����~��&��?�G&���x��9�O�X��J�,ݮ�3We�iD- ���>�c��ӿ��V��]���r��)䒢-b����{i]ֈ~��e���w�:?��؁����h��W(��M��Q���I����g�L�=��y���t��ꏤ�����9���'>i%^�-Ʀ�-.V.�.����;Z�6�wl �6op��~�}�y��gX\��[�����1BNg���U��!�j-�t�R7���BՓ�q�t�k[iSZ��	Dl�,�p�~5i��'6Q ��*8����Ζ�C�%�e|��S!ꊗ!��]n���Y�R�S��������o�x�w�����N<^i�ۣW���	/��n8���=8�;r<���Gi�P3*�<�_�\&0wlE�e�*q�_���L����F�T)�$��7ȧ�,�D���"���#BmH�z���<�T�q{>֢��S������!=n�ϖ����bv��H5m�r����p�+и�0��8�ޫ�t��*߈��S~l�L�������϶� kg�"��a2w��CJXRf&Ϩـ�V恈��n�K٪٣~�+�V|X��ݹ�Pk�pֵ����ѕ�|@�)ű���@d*R9q �ɝ;0��(\ڛ,¯���(�j�zt��|}��6�����Ic��h�O�v�ǀ�Hw�Y�
��;*�%$�5��y�8�k�q�d/��9ZM<Y~F�s�F���N���ׅz�q?_�ڶ�W*|�Y�:�a�G���^���mE; �TM+��o�r��6(E�L�	�UW(j��̈́�F�3ӰL� i��oV/�[v�ի'0���]5t�OU��k�#�eq�9�,��6��8����@@d�I�e������������b �����/�P�_�^@(�� ˸�X�U��p�ȋ�8�g�gO2q�³����g�����rϨ��|IAک#.�s*We�.�~6���qI�NRNAlx�bp�_'�uM��0����Ak���~ޱc������&�(m-+�i�L9�
��7ܠ,Mscry��o��jQ}�Q�XХ����a��-��x�g`�u:	�r��<!U��>��w�T6��1k:���|��ĥ
���];��Kw���a�ҵ��K T�$�q�q�9-�µ��I�o7%�M͖
���\YfǛ֤C:/d��oD軻hM�cH[��T��'^	jD*���Ke���lR��`F\�l�s=Nq�;'%��ʍ�gY�[粒�Q>
�ݝ�! ��ʄ��?P�� ����1���b#����c ��n۠Ӄ�n�����e�?Qx������`�׈`�.^]@�w�T�>��X�$�S�K�"��srN@����y�t�?V��b@��+���W ���}�F˪,�l~�g Z�<|h�v�7uY�V�g�X����{��9�^�sr�{6{3�x=�9o���"�1��ǉܯ�쾿�Da疒��%OI$r.s�$��ˆ~�^+�p�P	p�1�1{5�;���=�<���	�Е�t�Cy_��L��:���UĀ��a�h���a1�c@f�$?$�����3�*<�ɒ�\T� ��c� �}����1:cl��_0����:��`#=��U�<���,��JYT0E���e�C�w�y=�|y�dڿY��q��� +���8<ݔE��x���3���)S�!��}2�'��T�����"�ȧlF�{�&�;uTv�kX�颧^���"�鷎j>��El �#�����W8.D���^�*��: 4��Q�K�\!Z8��.:ՠ�j"��u����a�@�D4��
j*9Uo.�ql�>�`:��0n]l�L��� u�C��7�#u�@��R~\^_Aw���K7t�V���,�[4+�l&`{�ےJB�|��G�>6^�3j�X��q�R�LyQ���*KӬ���ɇ�9�\)G<Z�$�o`d읻(Wlj:��Ub��޾4�w�\��(Q*/�/�������I�9;��6�aZR~�Y �5R;���B��}~���r�o���N�uR �"�C��ƀ�4���+�b�۸�[G�M�I��}���G{n�j��|�� 'w�J<C=w��L��=�jF��Z�;����$����zXQ��Uw^��˄*�un�5�Rd��t�v�^�������^��
J���(���w4�<��nMysG��l�>o2I�����y�XK�D6g\B�$�Pf�d���濖����f
�o�����p�L�a��'A`���kD��7F�j�*����(ŭ����e=O@o[��Q���6��4&��3rRz}RX��v���U-��14Z]$p9Q�]��5��Z$��E�;T��kYyGB��B�Q㎊3�Y���p��kP����?�.�9m�.GD|@z�?�{@�\��+Ek��1W���+B�=�
�p�r}9
�p(��xc*�ՎJA^_�vGٝv�{��,Jx��}5�$�zg���u�a��Y�T�k?yC��h�bB�(�h)�l?�=s���hZb��_+���q���K�K�Ug|�-ǌY�y�v�4N<�-�K����NG}������S$�:_����7���ewdH�'��C�hA�b0:�3� ]�V�>F?�-_��/p �w�_����SR���� �l	���H�/N�v�Đ�㑝�6��c���N�A��2b���1c��pS�4�^2p�L�]߰i�,�Jn^�A����w=��S��Z��{zr��7�\���ȼ�H2ɟ���ԟ�� � ���2��C��B�[4_۸��2���EiB���LI�	&&	k>�E [�e%mZ�2�Z~��a&ݠ9Ig�|�����Q��g�#�KV�nU�O�/;�ą�A�Rld��<C�֪������d%��PEϥ����;�5"(:u����@�������wu��C�6�&R��QqپɷWՈ�G�V��x�=���+��8��U��I�+}�T�����}	|�В/�ksh�C6��Tr{�R�����e�~o�`ݢ^e�6̧�fq��0s�p�����i�6	9�C�d��
��|̨ ����ѐ�����ԠX�
�J��~' \���i�� ��,6H{��۴	��84����x0MW9[>��/ꟕ�nFo!��ak7�3.�(�`^̀~/{A!�玕�r%�=i-��8o
��l33��T�i홸��r�W�W.¡er��o�"�~�0Y�ϳ��	B��9�(4]��WL;.Cw6�O���:/����CMIg�����r�*G�����aUѭA`�T�q�$IW �7_�D�@$)�=)pڝ��X��!�l��k@y-��T�2�yY�?a��B�V�Ɣ���������N��}�r�^�(id}��
�W��c��k)��iŗ���=Hѧ�WO+?�Qj+�p%������E�k��.�$��H5-�^:�F�'(n�'B7�0ٶ	��H�U��Q����������Ԟ�ӯA(��5�m@Ԇ��%-(Ne&z����`C�Za8�Z��5D'��w�4w~#�)?e�&�:��XE���K��@=/y�_pK`�ͻ�0w�d�C�Z���Iٙ��+�yT�����9�P<6�
��`�l�'�$�bO0�&⏽��1V�}8��$��)+\P:fΜ�w�0��N���@������/��c �gF�p�]w��@ ��]���ea�z�-�ޝ���N<b�_Rr�@�'�PɥR6!�]�gK�yg�r]�N���ȝ�M��
�̣*�k'��>aZF��W���U\_T��i! 	���i�h�>�T}���*S�����n]r��97|�J{�2���ӗ;�oHK`��J�zʢ�r�&�0�%<���B;=��N�g�FEZ/K��쟥�j��P����O,�Wv�j�\�7�GeE~5Qjۄ#ׄ�������g�h�JWӵ��v ���A�)<>`;Q�q	��#�F�-֡�[3��ƋŌ�ƋgCA��� �kU�A�^��⥱6�ͅ=��Z���^�1fó_"9L�,+Tu�I��H�L(v��ܠf��c� R�Z8���k�*d}��q04��[F��Ɓ���q ��b�#�eW?`V!Iu�A�����hZ:��ۖJ��a#y��	�2�sG̭�s�����jHƲd�Z�3q��TN5f����jÁ2&� ���qᇙ�ʁ�o8�$�:ok '�h��J�|��ڪ�xW��`�_����	��*t����AY��եڛ�vaU(�cj�뼔B����$��Ç���.�ݷ��s�+I�>u���@��wd�Y�TQ�.��9�"A9S�^,�&�79*�Ӗ2 4A�ܐ����d{e���[2<���3�v b^#&��'w�<��Eo	q�~�������Q��:�,r�yF���x������ ��H$�q�ti�/Z��yx���KW9ǡ�^>L��2_9J��s]�� �_mP8kr�S:zxϾ8�V��h-}��v}�� wcm��
���)5�(�"��Kt�T�V~�{f���@�����!� ��/�����E���U'jR��$�8s]c��a�y��!#Y�e2��LF{!ύ�g���)�F���'�%D�B׮䷋�tӷt�S@<@�Ԭ����NvE��l�+�{���&�OLD<��o�����f��!n`��E/�y����\Oz����9�y(��D�Ydṷ�u>�\����Zn��5�1\��V�d	J��؋����;�_E��i�8��'s�w��j$�w)���w�ݱIR������3��]��=}54f+<Xܝ�ƺ�ߏ���dW*y�x&)��ф��^@�z,I	"��j|�^Ɇ��V?����	�\�9����� O�G2T���{�"����
bD�4���f�L�Z?-��q?���|"��i5���!$�x�K��ӧd�?<���th�=o����\ ����oӍ�Q��M�׸�odE�Ul�N��5RR׳rf<4
����~͗��0H�	���8M��.��gn�=],֧$�%�Ͽ�!��[��-֕�JL�t_��c�O��H�wx����#,�h��-�}T��P6�"]��/�l�U��iݯ_�c��'?�{3�h���м��z/klPP��*C�} ��K��]��(������,ə{<Q*3�KII��#��U6�ݘ0����2�B���2J$$��:8�x�Jp��)*<'S&z�l�����p��	=nC�_��W��:�f��6���E1U��"��"�<�#�e�x���t�n�"T'�4��c��B���*�m�~8����+>�ˌ�E�
L�_�����<�����m�5�j%l�cn����������MPd�U��y��dYxk3�6KG�#[�{Ͼ��A�any�%qa�b˗�cˠR �|��m���r"G�|w�:u�3Id�M�t��=	��%�6@,Y��?D^��R��&��X�u,�L��TY��N8�`ET*�h��R�s(=�H�چ���|�<Rb�Y{���c'&9*~������|�I`��1�e�O߅��aZ��a�|�&q-������-w�m����^�A��Q���Xt�]D�]jFa�y��ح��4�qj̃j|'P�S���u4M�T�"���v�6�D����m/{jKU��ҰL�9F ��Lwz��˒�F����+�j������V�!�Ċ:
��Ě�`�uZ��?{��
M{IL^��x�>~ �:��s�����F�6�k�����u��j�b"3M�h���K�G�I�λd��󝔷�t����ѽ.!Y$���3�@�,؋0�iu?YQҜ�}��h:���a9DyCW��F�A��4�$�-�Rl~\��=+>d���0�:��;s����	�����Z�3�<qEL�@�e涇���n񱲽ͻ���Z�E>���~�н2.((&��,�$�}��2�X8�=�`�@�������]B���|-�ߊ�\�@�N4]�,8l��2QV��ſ~%o��'�� �'��A+�<���ƒڗ��Z�^��Aǲ��������i0�w{�*��/R��plg���݀����� [�g�`�1r=�a��v^t扥x'����X+c���s7�%����V�fArm���L����4x��^�qR�����g�I��%B%���#R��w ����PZ�=�����M������>n?C �8E�xcs_@h�+��g���4��,9�����9J�L��C����pbm`��=��I� �Ӏ�U�z��'�>T��A�y��f��fVڎ�e���8��������.��[HCQ<���hdX%EL����Y����/��0uf?6�M���c^���|G�}x���pV�����`�"0���~ ���R/��%y1���|s	~:]?S*�z�Q�u"��x��I2��yҷ�϶fD��g��e�-lytO�4'[���4���&���l�Emr��hB�]��~���(�)�X��뺈��<�*��͢#�YX
��5'�m֠��-�DMFB��j�)\e���#��\��.�|�_�Er��J�^�c���|��	,���t�!�v6����	�&I�s«�k,�j�uy�<�����9��%p-�$$����[��!��#dq����h��r�e�����c�e�K��+���u/@YKQf�=n-�p�b�/sK�ձ��ѩJ�W>&K��p'��nks�Py��.Ĥľ&ӔO�L0��]S�"aWA.L�WrNo;	��)[iO�b4�ʜbv��/��L]rT���%HA{Jx�#o}c��~�������I��k��Zd�^�鐙�������'�p;4�s�T3�~��<����T���X�
�b�,���	�L;1v+�X���q�����2+g��Р��D��@�N���8�>�G �s#<��pы���FX�~W^��я7��]�NK�R����I�sI츯�1��#6�J3F���.�	1:f$N����A&-%�&X�S���)3(F��;�/mԷY��VH�9���\ax�y��{���k5��Rk�L���%���N�;�B��0
���cw�&��kqۚ�U����(+/�'Y�)r!�B��vy���w/0�C#9W+$�h������$"yi�$F/��J�����з����_
��^N�ٸp�SEH�@�c'��X��P�^H�ذ�����Tr��^yv/�
�r����>�ac|�n,�>�T�=�j��#��)$�$��\��B�� Yǭ���NF��T���r�DU� �D���_
I%^�\~͢�1>�V����@���/��S�Y5bN����u]�,�\5�%�@t�DyB�O�w]ue�z6��OD�!@����`�M�B������>����%�V܍c��L�t�
b]���T�W����ֆ�vwj�����[Ģ�S������1ó�@^��*o�pK�U��P�T`�ZՕu��0�L���A&'<��mQ��vע{�#�n4���"���)��W5�'��{���I<l���Q[S�tƖ? It�Ȁ��œ�;����)+���V���ޏ؈!�mIhc_3�(���'P����2y�І!���
G�,�~+����H2%ٙ=�Q�B�a�㿧���®F����w���?�J�LUt��Q����q.����*��I�������I���"MK.Ä�d"����AXbD�I�gz:8<��m�3ͨ�:��s�3�y�P� 0ʗ���y~��d��ܳ���.���I�����4&����"�4/�z�GT׿2/�}��e�;̑5�������d���s������Q=�]\Sr0C=;d�ȇ~���)�5=��@٦��C�$�N�D�o�RKi�ļȪ3�E,����5���w�M��X=;��9w�y���A�R�N����Ӫ��`1�9pN�]Z�a�fh3>��{�i�*���j
P��*ָ��#qY��A�⺛���g���>&���汦DwŤNYg�+ ��L�|*`�������Qf�)��C���t��Ц�J��#�u,w i���!�G��5>��J��;C�x��4�ʉ�kg	�s2�P���g��p򡑩��u.��s)�#B�Ĝ�\Ԁ�?�o7W@|��o���:+���T:?a?��N���'�O�c��� ���������GX#d��
�
�[��y�ȅ�@��C!�V��P|��K�}Ȉ�]Nb�`d��H�r����v����{�`Eo��S�J�b.CD���3�r��^�0�RW\�!)�_������q&����Z�� 9
=aE��ԓ�����w��Hٗ�l���
���f/��Ҍ�Y������W��y
,--ʲ�{���as��m|\d?��G���+D쉀G�k�(R��Ȗ~��ĉj�b��0�c��A�̈́��و�:&���9�?�Lh�*�z�`_Js3�8���۶/�����9�v�d�{qN�N&)�o5��Y��ՠn ����voƉr����!Ω[D�d@���*\��#�6Ɔ�a��>	]TR��n�jP����'�%6�asN}fD��n��D�G�|�;0D���=����nδ�����.���yI��G�~�L�[v<\����+�Iȸv��F��K(��֏���|?qF���2�w��9�}�%�a=�{P����e,� �͑�6��E�H�6������@��c�Р�����X�U+�,��u5��w�'G��p	i�L�ڐ�X��q�c�MZ�k�J�v��lh�7��<H���x����('z���-���,J�@��b�;�U"r-�v�z��n�ҿ������A���p�0JcP��(x:�&�o2�"̤)
���h���H
��ւ���R��l~�&^��O��J+kp� |Ã����"0�PP�3e�'���>)�C���>w��'�m+JmB	�l��غN��6W'���1�P?l:<�c:߿R`q��V���{������ي�1}�����Q$$I
v%��1�j��]�\9��Oq�N�E�,��l��.���q��Wi��L�q�B�*	CF��m��;�GΚ@�x[�7�?{�ig��Ղ�BC!ˀ+�v{g^���B��~z��;m��Vmk���5��>My�"*z3�k�~��M����1�n�ujw����0�黈t;����?7����WC�Y��H<�k�]d&��H�����6^��YiC���ū�EN�w�������~w�E������]��#�(�0��C�H�����Q�
w���8�vK�I�*ŀm��{<�����o�ŀ���(���f�z�������Q��c��@J���+.����冓<�6i�U�p��b��kP��5�aY���<�j�r�V m�sxNM�Ш�t}\�������fXԏc��J���Ws ��=�G��מqc���}�!wW���ٹ���W��U��N���J���x슨7�Js[t�=�V=�	?D8c<awס��C@��x6;�C���@96O���sǜtA�Ȣ�6s�Q�Sw�&;��dcw�^���&ږ�I%ώ$�� -�ϔ1�u�T����[1��12H�C:H�DB�1���e ��`M8�OZ���I�
���c�,H�Z:#mt~*ɽg�uE�fi�N�#�p�A͕I|r����]��z���s@top�|���DA��{���_���n�)q�)�g�Z��ѕ�����G� "��s�34}mh�q����y��M�RY	o�޷�2[��9��� ���a��f�ed�ڮ�a�L��A=0V6�v����2�(6��Z�Z �#p��4�uy)�w_B��_��1r����wx���q�m��L(�w�ƉA���?��M��i��<� ��z�C{^� iZ?��Kߧ0Q�j�E�T+��]#k2��B��m#ArMZ�88L��-7A"౑k�bHt��Ӭ��B�6a����s����5��]G����$�od�5����()�i�yY  �%�oߐ{S��U�	�&�8�ʳ�A$����;�_;��F���,������A��b%oe�7�q+�4�����iA����9�;�/���`�-e���=��4ȸ���Vj�pa��f>94mi,���C�8.��[���#�H������+�\1gE�i�qy_��btw�d�� q⭝X+�@�Z�2 �����t�%f��s	I|T��s:��l��yp�3���1$�i���;N���R��=m�u�Q)�J���mE]K�}�=S�Α�?�Q���_$�=3�}8��)�*�3����,3�|�2�>j��5 �՟�}��>�p�#]=�&���Ԇ���x �@L�GS��7sг��{��Yܨ��N�wյ��(v:�M�8߈,k��iƫ�ۡv�G�ɵ^גF���yۼX{4AN	�)XB���v��0�Q|�d�}��8�*�a%t9J��'�T�ѯ�nͅM{�]���3�|D{ �!�L09���R�M1�%�D,_G��e�o~�Xv8M}�ֽ�Z�Ҟcڜ*lw���"��dB�`�P��9w�߳�͗��t�Xv�:S@��^��G�$~d]4�(�{x�QY�ܸ�F~�i��n� iS�IqB��r��Q����m�=�<&Y�YZ�b�_�?]�v!��@�&J�Ǔ��n$�> xb����B����
5�B�}���Ǖ�Κ��iK_�����;���@i��蹸;�'L�'C� ����RS�NP��7��ڗ
%��yǤa� Xf�hz��ņ_@���7lYZ8ֿ=\f���"��5iH�#x̵'Td���{nm�n�8!o*4@/
�> &��v ���{��Y�/�� 
k»�"΀S̚�G��u=��u{!���Q���7�|(*^���]j�*�d���NL�݆�Uh�A�O �R�p��Ię���>�ΦX,"l����y�����专>`��0�)Q�Kħh�J��2���o���)#�f�<�i��
��,S�;�<����ؚ T�c<�FWG7���xǀ69��_�j8S �C��_X��\�>�;qu����+�F�vcخ��\/���R�p���a	Ev�S\0��
u���Q����i�7q�_WDu	�>��+|�}�����>�Y;]54Y>�f�8��!a�Q�@�k>�(�d8x��\��ݻ�uxo`�`,1P\�t�tb�:T6��A������ga�l�=�#�&��-D�ƛr�yw��%Տ� ��*/�O�R�L6�'�P�;�y�s{�9�=�/>d���Be�M�X�x"��h�����9�a9]?���O���ϋ���8	����se����)єI�B�?">���}�?B�ZjϾ�);�ۏ�8E�"���݄�#x�s��ǒ)J���N׳�h��,d��6�r��t��b���#�ē������M1n�ݟ���IsF��������T&�"����������[R���W�5����$P��s�Wj��$�b��%T���@���0��\�Y�vo0�Ì��:\����E/��΀[+���������I��T}�\7�Y�7ʨ�gyw��'|���_ZO[���	�꼋^��<�:2BkG�A1=A�MC��rX��>$���A��w�x{��U���Wn[��+��'Jؘ��7���������KB�@����K��U}��q�9����A��u�#Q4�	F�~lR<� ^I���%ǮƮ3T�{,(X���#	*ʰ�������ᓭ�V�Bq�m�*�ú���S�GߩóT�Ǣj5�F�Yʹ���_c�Sïn%�<�!�>�.n�">��?m�t¾�k󖘛k�zF����xb�*�K����3%���Ŝ��m����3S3��٠��R���'�|N�(�j2L�Ѧ��$ ZaaXƷT�y pz�	K�L���K� J(������V����{P�Sh	e�T@N��ޮ6YQ�1��G������p�sN�O>�wR''h�`)O�XUH���`�Br��~2(��i�pu�۫�#��	nU!h�T-��e�y�Z
��k��V����1c�z����*�n��uo8�۵�<����h �YąV$Y���:!)��h)�t,Vr
��C�B����z� RνQ\�r�� ��"H��14�w�2)��K�(���6jT6R�쟾_,T2�ȗ��85Cy^t�4���1x�t\�b���c�dD�L�ύ�䩃v�xXvCJ�E1��1{쮧�~�+}���^��u��3 ��A�i����{��W�{��Ĉ^���9).mv�ki���yy��/��ժ���*�?2c�Ou�_���b�.3�=����!�X��,�͇vE�پ��H�Ł���+9S��р�_;�!�db��/�d�|������95�w��½���[�o�%?CL���>\����[�b{Q�q��4�!��Q]s!�/yk4��cX�^�C����0��G�ǹU�m���Cܹ%g	��-��2'?�
? �A]��i��2��8/�������ڏvk�E��+�l�B_��F�9z�FHN)�h��-.
Z��X�8עM��
�ɣN�dL�*1�^���[�@��:���i.{���3����t�B9-�ϗb��,O����P���E�"#�w�P�t���,uR�K(���rZ)�Gp�斛/��.v	�)�w��ti�[8C���P\y{"t<�L�1{��jB�K����%���!$�{@_MٔouL�9�Cyl�N0�kr��IR����村O�Bv���!(�{��	ﲋ�W�,���9��!A�2}I�*w��~z?�^T6��iw�z2S
�x!Ha�U틹���\�Ӊ�w�djW�� ^cJ
N���#o$w�|�cj�H�uE���?v�= �Z���7ￋ�{���gn ��.L]R"�@��Cz�խzq��(@@.�g+�%��n:^wۗ�8�y�@[m��U���܃�����+9�����)T�X����c%��Ʋӗz�.�V�Z�)M2�|J|Ofo9�FEj�T�/X\w�eތj��g�;AH2�N	cx�ԝ��ցx?-���f(�O���U�Ŭ"��tG����(�x��,��%K�S�TU�91��R����;�ݒRm�ٻR��gxW%����w�`H����3����G�
�J��^[W�'��
��K�v�R;E�ϡ(�Y&9�d7�֎�����1]`f��3��lu+j����c4p�&.i����X���a �A8T?�{����U�)�^%�ŭds�7fd��IlD�	x��Ƭ���0� E�u.����G9@�ώ����L�N<�b��\?��(�7ʺ����c�m��0�]i\zHϯ�x3��Ib)k�,��j:��H��,�ʠ��C�v#����(9�*�Qb�z��j����9����ji��ƣ���5F�m'{�(T��b��f��q�
S+t��i�Ҙ1�v�S?HN�>���b���~��9�86�n�I��s~�/s�,�f���*;J��~��Ͳ����t������A�\���I����8C�g���(V���~���mY�Շb�v�Or6V��
dPC7��7:�[ڨ 3�H=�3�VI�V�=�����x�i�p��'1�k�����O��x;�\��8g^�vY�	O)��T��_-�D�s�N%n����/�&��v����T`��C7���M��Y�'d0��*a�&���J2�8��\�P�_Ź�����@��c��@������ߐ8��@��p��@��TG����7�Gp�H\��2�4�#A���7�~�vG4��������q%#V��X�ˠq��ֿ�����^��VQSJ���"c�a;<"���N�i�N�/������[�M���.A�C�b����\J�(]�U�y6����%�)�kp�><�����^��\��Ku��f*yE�b�M�h������GΤ�����Uw{sɧ!#��`;7x[LZ�QY�ڎ�*@�=nLyV.���-�ȇ�5\O�+� �tOSU��-�|����\an�5�$Rܛ�z�-
+��E���c��h�QtZ��Fz�Fl$L����!�3�_��O|5	�s��4s�A��y�U&W>��PF7 n�I|s�n�aڳ�c��U�qۿ�A�JJ���^2J2�$�e�S�`��C�6Yr��o��W�.g�5͞�;ϻn�&��V��h�4��#yAG�~Q��h�]��,�ܒ��� ,\M�&Y�r�����X?��P�3D�7��$�y�l��h
���/�Gj[BE�bc�)ҙ[Ox����m�:��s}5�}�u۩l�H|�Y%��Y]�^Ү�lp��x���e@�^ڕG���8��
S 9?+��b;9z/1!�Ÿ��>��e{JG��+r}�w�H��W��7����^�֊'XMz���i�*����F�ܢ j�X�y�K��5+pu-Xt4q";Ӽ/�_x�Y�4���&Qs��ˏ�|�����
��d��.�*�������$��i8��x�l-�H ��h�ְ��,�&�2���{����"vF�pA��&��ՠ�bH#�!�z��𱘨�a�9?���?�,�Қ/g�U�E��~�_� ��)��=�����|�}���cz���`ʙ/ �r+���b�pQv���:�[��K�$��k{����VN��߽�R�z�-�TnZ���q��X�Rt(��d^OETZ�_GMH2�ӂ��Nц�JHl;$=�k���� Ι4��@6�逸�CRlH��sW�dT.�ӁU�b�Z)��H�J{8J� �����1\���0�����
�Q���]R�2	��9�������X�=�. 8⦅7�S��xL"�����>����3�('��{U���Oդ�5��Q%�+��ʘK�?z`���:�����;�ﮧ�=��E�X��"{;K:Д��Ff@cFe�B����i���voІ*���8�l_�v��H�%���ܫ�N���z���:𭩿E��c�+�DeL�1�cÒ/$;���/eH���3��:��AVL�n�`��W��\W�p'knH[�$j��i�2�f[|��^پkǓy��� �RU�&^F����!��Gu���le��Q/�B�V� 5t�[^����t�Sjb_%ô����_�lٖiD6���u=m���c睨J��amȳF=�� z��p��B���d	���/<g
a���9+8��V7�͡��o�k9��?��Ͼdt� +��[�Et0��ad�U�"�1�$�Q�u�v>�D�:K�"Zm�z��3�9-�Ԑ+����Lun��������[`A�S�}?e.�^�
���8����!��w�H7�7(��c�m�i��?���2�HH��B��f�>�M����r�Ê]@�.`�ܗo蝊��-Ot�doml����&����&�^�z�
B�Ӟ�I����I��%!�|&� -q�d�u|��5��9=�jB;�4�jڹ��� �(~�|�f<wt��z;@2"��X�ʹDU��K��]���К�����M���e,N�#b�_
�|�xw�U9�[�#����d�a+�%�&�	��3i:�8Nustocm���*���s�b?�ӈİ�rA0`�qr��#%��s7��x
Z\��+�����n��Q�-k+�PJ�Ǫo���˂nn#��=�����pť�J���nÚW�`�Y��bgf撄s7��8g�H��am��h��(��:�?p9W:%]��3��3�<�G _2�'�M�V{�T��� �}oN8�#�l]UĻ��#S�ՙ�c0qt�\A��٦�o�X%5䍘]��9F�զ�X�S�?�7�V;��U�Gq��'3"�V.wrqT������ARP���R�����f����A��M�]V����JE�>�N>����μV*Q
���7O��$!l����U��$a-�g������"��%l{Ca�+�	j��;�DN�f�� ��k��紌��ø䂢Oa�FV\�nS)z�>����m���Μ/��������� ��j;u��c�]H�2Qx�T�2Z�j�4�+�8��Z�s@\�H��Z����㚜���ndbۻ$�����B��kP�JU�?Da����	3=
(�kܗL?*F��XF5ފ"PJ���-
F1�	uĢ���I�]�[3�o�����c1��D:�L���#� : ��]��W����u�s��p>PGك�7D�_���!�O�̉�<��B�U�=g�rj� x��K���[GY6��^�o��e�LRb�r4���tO��G�`P�0�~ೱ7t��˫�K��~�d�~����5��G�r8?�!�7�(��L��(V�TM{���*Q2�mű�.��主��+_���Y�,�1��9��r���X�N��l�of�T���9�����av� ���U�7�n�̬��<7������IB��&s�sZNcv��E�΁v���=,���W��c�]�� ��J�,�i�"@����]�{��+~��CG��VpQ
}f���a��yP��Rv���zt�T+.B@��+�U!:��9��!��|�u���d���`�zj�2)�×����y��<�ׇsghzYT�C���V�e^Jd1�O[˻\���Gw�bs&.7�ȸ��vG~qq�n��\��ܨ$��~�N�z���IVc�4U����X��0۾�ͬ-JJĐX�N)Q�d��k�b5(�J3/�<�oW\����s?�$E��H���o����%9n�e���)k����'�&R��3�`%�����!C(��T�τ.g�;��q�]hH���jFl�����{U��� 9���p���>��I|�^gO�H��T�psV4�����������`��v�K����03̰Q�	)~]ʤި��p��W>�?�=�LQ�OC9	?U����k�jb6X�$�'2�2|�e+�?��x3��\����=X�XD����b��rz�;h�E,���+M���*'��u����&[����ëN/�TX���j�)FĹ��Q���j�W��6������T��]�^Y��pkǗ>/W*����סTO�0*�x�d��O�
0���K� ;[`=7/_��ɶ�t��e<�iɻ�;���.�pY'��e8v��s<-�]��������b"nA�jk��J���["�1Ӽ[�� �yw��K��x{�@�@f'�<�~�vĀ+*]:l�v����g!�-��"�3A�>@�&�m�x퓞 :Ҵ�����������&���	n�ͬ��[3�O��$@7��BPQ�w(�AH�6Z)Kv�����,���>W_n
y�B����bA�9�����m�,ܼ:��}�*��6�o�hİ.���yR{R�\�[a�Na��$n��Tg���'�*��^�O� e��� ��u�ۏ�숟�N��'�;i���7����Y�!��� �C�e倄?���gj���S)�M+�N�ӊ�*����ǇK]����ׯ�)wEĖ�����	T-}� #��ft��~���PD�e�HB�	Ve�����"��z���T�H(���U�|�����tS���W��>�(c��ï���ŷ��S�$r�r��F]?����Jb�X|\NS�px�<f0����"���+1��� U����f[,S��O6��ƹ�o�f%xviBjLI��t
���J��݁��M�/]�c8�ޟJ�YF]ëS��U�u\G���7�Nש����;2۰U�=����y��Y���8�>>����e�2>5ʿdc�ذ&"!� �d{خ�U����|ؚs���w�	u'�A������e�}��]wE���ɠ&|��(�*9��!%Q�sg��<zs��Dg���{9���ڀL>�L\73"���f����g���}f����~���#�u�*�Nw"�m!�g�^�.E�<y�����79��+o�Y H��U��Nw?��p��������K�^�:�R��:<�z�Pޑ��ߪ�n��|<bzo�hW�9߆�CI_���?v}���ã�Ls��r3������w�� }@@���b��P������x��UC�F.a�����8�����;=3����=ky5�)����C�"���Z;�G��U;����1~}:�̵��?�5�� ��x��p�(0�l��X���Nh��M���µ߂�O�PͻZ���6��<�@7a�i˖��%]�(�-56Y(�-�H�i��8�=�+�2����s�M�	U��d�;���p��k'A��8�>�:�x����T��W71g�h�gBA5�ާȾ/���:��@�h����p��5~�Fp{�r���S���MdB��":i8���>����\�,�����k@ ��C2�S��F\D� �0{sR�(lq{O����m��\�z�?bI����-�{����G/U0�1��;�����Xx���3�5��4���:����y;$�I��V��W�f��������A���J�9OL�3U�~��������|A�S/s:�����ɎK��9~�.2t���F�%:g�?�\p
ꞌ�Ȉ���`���&j��H�����^�-K,�I�>/���d�*��x��^Qp�0���4�"*0�;�kL'����6)�,8��mƲ��9��+|�"�wxo�ꦞUK�Xz4������TG��6�<,Fc��f�T$-$��z�� 9o:��&v�nѴX��ۙ�<[I�eH,S?�bA�o�9w��(�����A���4}\C��5�!���N�3�ѡ�.���gG��	�-4�N6�D��ފ���\��=·n��5�<B9����1�2\�������g�@A��Q��@H�*��Q�T�5%�	���
�W����M�ד(6i��[Ƽf�9ɜ�}y��^YI���l�����(�ў�0gu�����i��E�	=J+�=�N��Ҙ*�m�_P��_tr�ƦѠ	OvG��p�/eM��X��!Y7ʲ���1.;�j����{S��ܫ��ZY�OB�	K������r�^�(�D�	'(��)��Q�fY�*kp
"����t`����6Y�#LzϗDo�����F-��
��	�B�������V�5�~�5�hab��������l�oԂB3�AZTk���c�r��My5�X�+!��/��s=%>�Q#/`�,jXG�r@-��>�}/=~� �Q�Ipa�]e��B��.9&@1m��#A�9��K����,h�I	u���8l72A�Prb]wh��o���,ꂾ^^��V�Cq�2V�Ȃ�ҁ�4L��9�-O��}W�� �&y��^8�^����zZ���zB4� z{c ��vi�O��6����K)�Dd9�Ƴ��5���R��x�.�!��c6n�@�6�AX�I��HŚ�b"��έ�#�rq�N�yN&��P�$��wD�G���W����U�����g׍��ut� 1��0�5JT^�Zv������SAOǢ���ƕy]��m��9W���2g��Ux�������5V�#�?c���.�͠K�
�� h����TW�V�AK������Al��"��P �~��)'1�_��7{+�a+�3s�s�d��啰��fmdO�E�L�1�΃�^f7�� �zP�M�νLޙJH9ھ�+#���3\�{e�J�I�$��3E��EDa�!�Et�<G.�`��i�uBh%Je�ճrd�q�g��7��B��R��!���c��� �:Ba���L����#a$13Q�[�k���og��7H=j�s���6�S��f]�>���h�e?�ݤ'��Eȸ��"��@��^�B��9���0;�����e�$�ޢ�C � ���h�J��=�`��O{���1��!7��+5���y��3�ዬ��8�,�!�8;�dE���u9M�5�-h���~���6�}R���;��52ay��]�
ӌ���EFe_TG"��[a�שOG=�z���{\%�Z�ԓ��Ѥ)���l5��#惓%:6{fg���«	�(9j��s4�~��r���N�P���}�k�BCc���P`7���c�<����1.�//� F�����'_�b}ŲI�y��^�a� t��;�5b�����|w`���^������v~�����Ա��C�	������e��y�z�+��9�!�ߧ�d��mp�^��:W���O���� @�k���"4�'��'�,f$	����Ƽ],�%��]�\��	������fޚڝ/��Ї��@`
�{^��S��Q�^Q&3|�$Iİ�=����GSm�o�@¬�_6g�h� V/j�Ξ[ �
HP�(�W�K��澜�$wNS�Y������2#Ӂ�h���\�q
�N��u2iC���:�msA�^$�Q���qCgC@���l���~��Uar��x!˽7�||�s�]����$�r}��H���tf1���5�w�(�@Bb��*���Z/�(&2/v�P�+nG5��6C�={|"�¶���,t[�*���ؽ���O�"�×:��Y��#�`�'0;iǄ���}'b����Qˀ<�uG� ��0����@>��(c/u���Z�^ފί8��_w�kq Gk�M ����Z]!-��h���e�����.h��"�mL���>r.(&��Ԩ/�v�ӹ(������D)޷�$x���%����:�E��H��Pa�6�XE�Z� -~�ς7��,W�]E�����ǻ����L��"��L|/�L��g�3����%k-�LQS�?K&��p��_��+@��Zm�C[q�2һ��J���?��%���-2'f�
M Ģ� �u��0���UM\<G���x��}+f�aHS��֙/����~� ?L"�1��o�s4f�3�zlŜ��31��;-��h���E���,-���u�g��^�oNY�rf���G�h�Ab,��)#�8�K���	��m��Nᆃ������(��Ao�x�<M�}i�r��q^�����*�d�c�>���m���9nۋf��> پ��q�{����0+���ك���-7��1'�����4N=�	K���wx��j=	�@�7Ƶ.���,�A�M:Yy�����w�αi<�⃥��P�F����Q�5�zb\�p?Xے�BCK	,��;� ��U, ���6d�*��+mY��{��A�~eR�MWbP7�Rez�-��ѫ̤��R�R&��uR�+����z�C�Zk�V"B����fxm"(A#���[_k�����P��{���y��^��"�/��a|aζ�8?���=�[]f�?�ٻ
]a^�t�&*sy�{�������O����>�ԺÈa+g�ѕ�yh}W�BlJ�9̪�4=����"���{�%������B�[�bn�S6��f��
�r�<�R��c�?�ݲ�mX���q7:������;;I�S�;�.���d^�4&��� ��~�͚���s�l~��|1.��D�z���P�TG��dH����p�|�#t.���M���m�m���ȶ��F�0$lk9i0:J��+�FW�,�����h�:��\Ю��.{d+�墪�P�߅C�F�3�s���?q�L�$t�\��zT_ ;�3�ű��4�����aEj����h,w�=��k���(r�w>���/0>�J��7���!�W�%U1`�ɲ�&�ex�6Ľ�~�\���z�`O.���N��� ;!��[����`�|<;m>N=VW��\�|�m/y�3RFa�~�����!.F�y��=�����P�]�hÚ�&��|}_&q���x�	�`e��30�	N ��oޱ(�����`�R��N��
ڈ����H���y�5M1?8pGV�b�:T��B�kj𯕢��(�9R{Z���ƻ4��i�P�� ���|�Aƛ.4�����6%Lv�h����(�[}�E�P��E>�X��$c_w�>b�֜˻j%A�"����6Zv��`qH�e�e,�-��:��k�v6DTy9xD���6�R(�J��fd�6޽�<���<矾�'��bg��1){����
���=-����B>�������ٴ���>�vuMS:����]U�w�Ivɳ��g:�ia���� ,>��rB[�V6�Բd���E��7��8��r��5.�a[������|�Q{P��ȣҼWi3�j�{q�S�fH=6���(�B�$�����S�左�{_o��l�EmF/��o���W��:�t�/ׯT�V^��C~�Vj��� p-�dbW.r��,�
��#�oGX�|�����J��%�;�W*���^�8x��E�>2����L%o�I�D�ρ����Q��<��g��pI���]�y�ބ�LCc�QϤ�X��~��<��r�F�2���QA�S�粹����Gz�ۉ���4�ÆJ?�E�ַ ��g=�k���9[{#�`��b
1N1zX{	�B�R�W��X+Jz���f*��V��9H_+��r3E;��>��z�N������|2���V���2d��ҏO�e�e#�XX2�� �BC���k�4��k�d<��J�,�i�Y5�t�I,��q��l�ň�h)�{����c��'�X��6���(_������л?������^�;�E��[Ep�pX��23r��dIA�������#,���k���VO�x�ᢂ����d��8�.��L �Z��5j�_s栓d/�����A��AĤZ�Z�D�"yC�t����Ro��Ԕ_o�q��|&�:7�N��C�L)�ϯ�|��#ߴI���cR����(�g���"��|y*����t���S��pc�q�^~�f���#�����*6��:�d2����U�Vh������O6�D�E,�Q���O�Wd�n�<hx�¤oI����2��E^j�TF�ϼ߀��SɎY���&���ugk?����,���`Zr��Ao�Ħ�i��bV5�<ט���\ڔ'7�N
���E�_R* >ؖ<�T<�Nbв7�I���E������-���}�x��M��Ewb�w���;�.���5@.�N+>L��<XB�"M`$���hzw@H�a�![�6�rn
����ڎXA߂��ӫ�EV��!&V�,|9HM*�����G�
�0�ɳ���B<��*7j����XL)���E��r/�QF�
�f�^��[�e�U��8f4]8FI1�%�َ�g�M-Y�Q�5�N������s���.�V)V݆�W�SV�LP+2�RZ= D��_K]�ŵ��ȇHLd^�*/�Mmu�m���~d�:� ����/���e�Yx
�AS[G�4��0u垺�ɕ.Ap�k���E�f���:�
U�^t�t:�t�����J ���\�԰�v9��^D��[ڙ|B�__9;��y��J�N]0�"�6P��7KIQnc-JB1>�uת��h#�>�e-$���t �_���y;��ؾI�Z��#䶲Nϗ2���驣�=���}�7�yě��7Q��B��(A�D���´4��t���"y�:c���[x�*½��ְz<����5�U<��p�d_'X�B�XF�Z�;~P����]�yn�%̳����BTi�%M�w�섡/ ��{؎`��E�9�FY��*P2-���V4�"Οa�Wc�-�����J��fF������Ǻ�_@�)F�?��}sp��<G�����8Z��ċ���*��"E3�bB�]Xr���M��bm�����U�ۜ�М>=Y��������Ҁ�tGy?�nOn�|�zE�\I��z�מr�#hW(J�:��(����¡�S��r�����*�w��vȘΕk���]X
Ԗ��O�uP�
��HxwG���D��%���$��^��Ӛ�y
�ǩ&)�j3�C�(X���x/���)B��<��=`y'0]u��ĮS��Q �2�1�jʃ�WU���M$8n��Zz5+�+߁픫**"C�u �҂u���)ћ�� $kLvt^,E��L1STY�R�&���S�B"r��Ԭ�G镚 Q�}K��TT�*@�O�C�ӽ`���8H��R�����n��dCA�'��R�!/���݆$����NE�t��_V2Ѭ��2ha���m^{�{1Ѣiո;~�#�T�����;(v#���>�]�>G9=j�۴]���U����|��_-�?�li�ǩ����n��%�c�^�.-�ϖ��n���(�V�q!�~	+H�ș�{_��T�cz�ɤ2�ٳS����}0��NZ��w1��A�*0꾜mOyM�?O�'��w��S�WFz�J��E��	�i��_�#5�S��Fa�m53����[|��qSs2;� �Q�fmjǤ�U�V́�]���}U�n�ƣ�O��gR5�@h=�j<ED��^��"'��*�-e*�����'�Ɨ
�3�X��ޡ�:生yo$E�f�Th2A�4�4^jFL'�$ȇ���!�P{�Щ��(���t�Y�9	��^bn�;��=�����[�� ob\����bo�/g�wťc�.F��ρiWm����|�Q�<�r!�4Ч� -^���ab�7�T��}�����ό�/��7�X���5���!�[`*A�;���rm���q_sD��"�v$�j�ZZg�b���^�{��|(q#5K�i��͓'�{��]�3X��}x2���F��L��9sQ�<�fZ���B�;O?��!����)���_�G���>�i���/����+t#/�v&� D�`�Sx�^���Bzi�������iX��xъ�!��f���Y�;����M��	�����c��k.&m5��'m�%��bn��E>=���ﮜ��r�#A�\M��1ev�%l�rE�U3�P;������lNee��w�	&�����Z,�a�nowQFlV��� ���:a�?.���.���>G���&�x�_>�`��<�?Z@Y�@cV�q�hmO�C���,7ly��"{)0���1q��Re��Ω� Ô�o�2,UMv�.��W\P��C�)�3|7E��TJ�t��z8�aQ/҉o���s"��8�$��=�W��;_���*�f/n��ANm+[3�h��jhjp��][�>ew|�8$9�j:��S����!z���il�L�A�t��/��T3��u��<��-7X�r����w ���M�4MaxY9�c,��$�o�%{��P6��'Ȅ�e�n�|�[���g������헦���B����+�m��JxG��˽Y��|a*)�Z��}��V�t|�O��S`��%���o8�)]ʒb�@y1ܘ���;t�s���`�U=-��8ؗ�D;�� 	�s͵R(���7h�',���& v��o}��_�*���4mn��L
��i���0�\�m��\�K��.g
�~{��d@�
������D�C@�!sc�' ��M�:fF*r���aǾ&<%��@�8�☬���U�~��~;�p#E�;fJ�^�-+��^�;�F�bB����K]���:�)�V�m�8�u�6F�N|8����V)8��^��A! \ࣕ ��6ٱ@��I���Wޱ�ð t<[kaJ��'ϱ�϶ ��r�ь�*�>I��.�5P�|��Q������'K��<-?��w��X/� �B��
zţ�G&�A�|��JYD��:��9`���`>K旡��Y��F�����=�.|:C�gS!���|,��

ʀ8��z=K�3~vs����1n���2a��IT�ի-����[FoT��F�l���dz����I���?��9F�˹-w��V�FW�33N�;/s<����.�j&j��!�.I�ꨐ���g� ���S(ho��Ak��:�vY�r�� ��>���S���i�,���D ��wv���ڋ����a�:i�z���Y;�0��¸5��F� ;'d"�U�+[�w�����B���"+2�TP¢�'p���H�ב۱�P�͒�y���2m���V@�y��R�6z���$Pfg\��V1����ǖ�,���`;��"t��R��a@a@9:�,�]ar�x�?�+�j�n��ཚ��1��ܿA�N1��p��ec^�]��a���� ����a���p��F���� �j�X��yC>�\-��+]�9}��eI2 �A�fZ�J�QL脐ٳC���n��T�ڌi�����p0���<[݉�#��YH^�W,�y!��\�����z-�n�:>��c0�rօ*;+�*�/�ˑ�9օ)��a����np�Pо5((t�]�t���SݒV�l{_E��:���<�R���k0h��*�O�~;Lw��N'�t�pZ��?��h����_�ǞC�6.�e��T΄vg�����J�fۙX��H�,0�l_i�u������),����%��Lc��+ȱ�G�U���b!�)����;a#���x=c�У^V�9������A
y�ӜLyOP�����m��2 �<��w�1ס=#�ObBG�&����+�gH�Saot�b�3��&�:)=p�"'K�U�#�=��4k�)E!��$b��mU���m���������cj	�by%��I�oĈ5�Å��a7���ex�aL\Ave><�kN$	�G<D�A�~��g]BҐ-��)X�¼eob7!��{��K�T��yJ��6��]��#/&�'�d�̿�
=W�/�jX+�?A��],[��?�j���>�(H�	t�?U�j�.c�R-�_j����B��s�i�GҀ-�➒ƴ(_�1�-p�{Aj��1��P)V�8DR<�������'�R��j'r��O �{��$^�j��v���%q�\��A:�[���&�0�&6FnC��rsG����-���&ݢ�)�����S'�X�WeŹ����ۣ���q�@ l:V�D�7�헰�aR�L��}�hЩ8�l�|x�RhO���Y�z]-)������<�	�u� qd"�K����O�{~���h��N/Ы�EQU�Z+߳���K껐��}���흗�;G�MN�
T����I#��V�K}��n�{��u���Sa`�j1��;1rxRU�~��TcHz�f����h%�	��xV+mQ���x���:ѐ=��Lj�g4,�`u���� ky�֍w4��6V �`����iS�~�JCLmdt��_��@Aʫ�.� k���hͦ�8).�&��#Lqܸ��Ġj�
_��Z`���t,E���|�r'���,�o�d��V
�&N�;f�	r@�4�`�kZ�U�T���O9�����$��4�,��O��3�~�{�1pBx��g���@\"�_w�89��U�C����&��4��q�)�̏x:�#7�eU��8�Q���l]�?\{����.�ո��K��9g��y�
*ezq0��m�kʎ�m����ޮ��¥P�kt*�X���V�����W����a�[9=��u�_�RVji������;���u<e�O�˵�|�0�"Y#�=�� z2A3b��2�cf>����f���8LZ_$Q0蕔=l�'��2{��]ՐX>�p����"b8����p	�8��4=g�}����
����.�]t����c>�4<X�H:������e	���)#����5��%��=�APzx���|ʕ]��ރ�Q���&�LQ��S�8��a��)�N�/p�E��#�����`l{ܡF���,St]����i���Q�U�2�e&ʹ.Z�T���@?~�	���:�f��X�̬�w�����_����.9�К�ʵ��v��ZP ��!f�n�t�1��O�P��fO!��M1�)�r�BEҮ:��,.��\݄Q&*�6���:����Q�`p������s	�x����7?�#p�I&���>��;��N���r���)l�����p'��2]��Ҧ˴X�5�i+.�ᄙ�X�
�aAD;��'[�d.��li�F'���B,�Y"`�D�K=�|��@���@�����&0>��F�8,���?���@.;H����7J��a�p�m�3�~�g����G����A��8�\�w����W	u՜><��C����"����=��~n�K$W�,IpNƖ���Zp�l�����MQ�%mG#\�;<�h��]���7�N'r,�tT
R�9�lH�j���+"�T�ړ��d�;�,Ը��o4C�Y� Ux��`AZjI�f˃���X홬�?�����{�=�R�cN;�~��%�x��ݶHj���_��3G�1���w�X�d78��J���^�z��j�f��6U�ckxV�J�*��Vq��&k��Z�ެ.MC���sEԘ���nS�Ȋ�����Ce��0?�;�����Մ��zf��L�K>�0v��6�e��Gw���1�sR�,���s�t��9��m��8XY�6dD�t�8 `)h�C��ܚgl�V���+
�+�*�a�o�
HE���ڑ9���޲�o޽҅�;�z�L;v�a�Hj)�#P�ﵤ��r�s���c'��o�4c>,� 0��1]Ń���<M�R�I(�͗Ĉg�0u7�4V�5N��O�uh7�*~B��w�F��1� ����gs+�R���}]ԃ�{�̦�X/6(�s2KN O�,�.��[ot{� ��޻�*��g���˼�<8%�n����{�^�l���R�E�[�$��ÎIB�����#�ߖ0$�<?=lʓƞH6�de|�߾ �z1d��`��'�&�p�����3d�o�#���D����S#����ه�)��Z�I��b�%�U�Q�LŇ�t�	�_��wG彔{����?�Җ���˖ʟ
Lg�I���kcу)[wr�sO�;f�a���1�[~j��X{8�Jh��6�qk�O��0@2��
�)`n����2��YT*I�R�}�#.1����z'`*yY�ˬ�������vy���e�ۃ�Roo�q���z0��#0��1ԃ�����w�9���0�3��Dö�/]˯��xU����QH��#�1\ƛ��MW��t���|c�(��M������a�/[�e,0l4P�$��I��u�=X�Ck�N^��Z��B^/�J(t��~XMb��J���p���mI�5�U	���4����������GH��q6��R�/Vl�N q���{JWJU��۩E�(2�؋qsV�;X�S0�A��wR��-���G�v|=���]���8$��^�G���de���x϶���N��m�j�y��/<��΂<�D�sgǊW���>K������{��n�\v���4��`���'2=�$}��}b������%W�3�eE�U���m�^��=[��+X
�+�_�"iս���{e�z��C�,�P�)U{�<�JJLcW�"*n���'�
OşH{+����s)ФI�u���r%w֪8x85f}�z0���UK�����&d��q,͖���d�ӲZt������.#CsV1������PN�`����Y��&f��P�$G6Ӝ�/ԁ���Z����س����dK��r
B�~���	���5:�:��£l>b'Rv}(ᗉ%�c�4�JI�B/�,f%N�PmWujE�@�෕FP��rQ�sV����$��k�O@<Ӂ�߶"�A�K�U#/r^(nY�FWK�-n<$�Bw����L�+���{�g�&�>�6U�BDQǽ�������Onoɤʓ��F��zg���.�=�~����Գ��j����:���
����}Z�˦D�\u�&���������v������'�������*��.y��l���6�&Ee"#�[���(��	�}�P,�Pkl�ŠP���:xΫ@.�,����Ƨ�ŷ��>��dU~n<<�K*���+�K�B��Ug��:lR�����jޙTI|~�]��ז�_�˵������+���+0*��H�V	��UXD�{��x���mެ�:��|جv�l��W�z�GѺS���ƯkS�%�����Y�ȥl��w�����h�|�zKu�S��?��`>`��o�wĻ{626�Zܹ-�!�Z�Ī��a,�K3"����hD<mUD�����~$�U�`1�R?0���My�����
�y!�.�c��|�ؽ�\���kC��R���q�]|� ���s���Ng��}n�>w��i�y߱NVghĴ�k�C��	�s�pe�L{K\�-ꙏ~��O#���M�!'>k�rJDYu�;�4�BEޓ
�M��#z���QP�k���i����g��<;�'vER��Ǽ��k��d��۩��A������ы�d?V!@B+�W�?�ui�b��}H���K=�"be��s���K#ȣCe~�_a,����GɈ�x�{�ϣ�C�fB�̏�88u�Vj�tC�j������fxTKMߗ�Z��*��O��­˘���\fZQdB��&��=�aH e[{0�Tw^�WRY �lfZ��g ����1У�/����*�%�B<S��$�U`�3���n@1Q��г��:���}�l��Kv���3�1���hU���"� �Qgs@#�C��(�A'��������`B�ahAL����v�֡~�#J��x���j9;��y[��c?|� ����X��ǭ�,�����6h��nF�Z��u�����n��p+�)�?{hKPn�\=�E���glǶ���e��� 5�	���=�گ����܁3`7PuI��J�1;ޘ��0'͊p8�tN.b���t94�#9��K��f$��w���d�wHeVx���S��j6�Le;Cd
�Zj��8�B)�t��$J�ܚ�}����:�m�)~Ш*܂�s���B2XHRcqm�0w�0X����g�LY+��F��O9��`�Do/�g�]י[�
��!Ė��6Nc����bn~~��Lr�Y	���4�d"�t��"�S�Z=��d���!N<�d��� &Ծf�Ը��]�Z� ��4h���J�TmD�� �ݨm82ؠ��*r���̖�}��J 7���� T�_�3/�^���_#�p�D��E*�I�Tafa�}�)#���"�ǝ�P���u�(�~h�n܌��
���r (]��O1��������y3��7�j��Qr�Q��؋��w�&*��= �����O� ���b�)g�_��J����߀j�w��	��Śz!�������d�&��Z,���u�s�C���3ο�;�Q�%�oÔ2[4��p��oʫV��"T���̏�"��!h�"����L�	F.�M�C���-��͙M-3�Թ�t��r���JI���c�>*����`^����^��u�X�ЄЏ��B�����n����I��Y�g8�.��@��������}�0��Stv0��CH����6���*���7�s�f�Td+~5!X�IL8��>���Ӌ�lՈP	��ƌW)8��a���+�&�nE�a�����e(�z"u�;a�g���l��~���C��];����= I������!r��t��E�@�kw�@Y0v*���e﷽�.�m��Օ���*�:r?�P����Z�WpІ�8���=;�����<Y[�>���wTK�U� �!s��?�ްy��-��n�L��(�L;!�d��,{Ǵ�4�υn�u_��9]H�yXe)�i�*<��L�(�g!��>���b;���>�5zëy	C`J'z'�;0q�M(�"�����^ͼ�q�/�m�l��(9�YS���K��c���D�*�gJ��@�o�h�/��i���!2��W�y��4>��/�&_�6|��>/�t��[>�&����ʌSQ��f}.&�lq���ʽ�!�u�Z}C��
I�0��g����N�n(b\��)[����5�d��!����\B���,<�d:c�-[[�~�	g�*Vu�5!1.H�<	��_�&�g����^�	�t�ōe'O��j&CVY�#v�mOj�s�� �C%�8��'��PI���ɥTv7N���Le���'wl8�N���0[��=�x��e�yEV�]�����U��	��ڊ6��q����t��	�b<�g���,�A�.W�3@�}�ֺ��:{Ht�$�	c�%�X�%�_��z��tT�Q9��=�#����LF�x��#�D��y�<c�)��m�._���������=�o~�P�W��.4.�=پu�cD��
RWYS���-Kѳ��e��}Y��V��ڳ������yz�RzȘ+̤����Y�R:Ve7�O�vjE��n�g1�|"�2�k�M~{���
=�ɂ{��l7N����N���� ��˔�p�1�b"�_m�S�H�x"����a�Vn�ʝe���n�$���a~&�?�1�%�@��F!]l$t��5����R7�)����X��A׀����%�&�+�ʵ�/��b g���1X�0q
'��5����K�M�	E�-x{T�4^�̂W<�'Eg�sK�d�_4P���##LJoUĿ1�7���C��x,M3H-����SǫEk��x�_픬]~)��p��%�K�mD�s���f|���?PO�(���4yU�b�H�3=A�Fd�9m����L���3���ς!�����m w�lތ�]|S )���ÿ�&������Ar`*�IkQ;�C߭�e>���S �{`�Ԡ�(6� {ΜV��H�B]�O��֒�5��C���'�+3�*#"��ȩE?B��%�/4�}g$��gJ���Z�<Xć��AP��e28D$-~�}��G����pIw�OV[m�Ph?��C��3zY����C-T��ԯ�E;����C�2A��+�ݗ�-��9<�9�}���֦2���V�`������${\���a��7�v��A�?�_նG$�Ϟ�:�J4(�4g���k�T�.�k8�����y)/��4�p��Pd��^��)\ރ��G}���������>���2��5;��`�����H8��p������X�CIm���߉Zn_bW�?I\�{�%we�Jb8�5>���`��+R��� �Z� �A�jxq��)�<��4���g��']��.=���T9Z�`G��Z5�K�X�H~>���%�ɾ 4Q��'x��F����p-���4���TFO�۔^S��H�Ct�*wc��n
q�ԛ@4�����Ex4g<H���&�~�?������T�3Ϲ/p��%�OML0p��<��Q���ؖ��>Y�W��B������B���2V��;�m�����i� Ĕ�������� �wA���6�h�X�ۍ�,h�w�X����&���o�@�$�(����Y桄�S����=�2&�Q�~���+�� �ȸWU��
W,��$��X���d.�>��m0'\$��W"bI~����Ir�O�;�9���1{PRR�/�Y(�dR[���U�vV��xP������XRZ��p�~JH&�ѥ�V�~�+�i�8��ʮ�gI����D�)!Yh�) �:����?���IUVq����n$;^���ML�q�l����M?K>�I��͎`o�� dv�ңOƉ��k�m��z��-�uj���aD�{Y�TM���M~�'Z�/ml���� dh�����l��]2������.�ӂ#F�����eH�9o�
v	1�89��YG�;�d�K�=��}H6����j�w���X`�}
fe�<���!��*�7z���������"E[L���s�<f,�Ap������8�]�[�T�|�6yƴ�Kgv�֗��y8��̀v��B��lP(/�4dgix�/Q���ͬ��h(.�ɕ��?X�6Q���2R���k��*�7^�gx�w{.k]/�M��D�dz�C�c�A�<ə(`�B�?z[Ew;ҧ���s�Q�*��Z�ӓmdGͅ;b��u��ci�S�Q���O�w�3� �%����髅��b�\F'j(�����z��B�Q�h�I��OD�j�[�֓��"��-R#��^�f�~?=H"�k^,�*� Ǧm��zeh
�~�$7�N��~�tX<���j8�&hӱ�4��sB'v�Bb�s̯'� �}���	Qrh�C�,0�O��;�S���)�D7�+N,`'ߗ�.��?�LtG��{5 W�+U)��D�7f= �wkB�������
�ai������R��]I�����xk¼��t���;uY>�L~>��L����q�:�FGiޱ���Y�S�4�l�\��Z�>�Լ����)��,:�����KQ�(����x~��;��QF�2�^o=(���D�hK��U���Y��*��:�X�մ]�ls�hb ��B�h�Eբ�,���z�" ��\$�i⊋������lA_Y�֌%�����`�`ǗlYP���k6��Ц+��؏!Om&�f���H�h�.�U���[�4�-�`	Z���
2c/k�Q��t�q1/�_g��͏��Մp��O�\�NЄ�|ç�iK&
�#�xx��񴉬ᚷ���]�вA)T\ Χ��d�3J�)x�6�Gv��G$��5��:0#�fn��#�kϻ	��]=�s�$��9-�0�� I���Ug6	�����N��j����)0<�=�2m��DA�ي���{-P(b���f8�4���o��ga�	`������Q/m�([{�Nl�1[�]��U<Q8�o��G���y)A���z~��N2;T��mj����^a����B��O�"<1��r�8a���t1dZ�!8�#��S��2��U��: ��W�u�5�2Os�	�Cv����EFHmU4Z��E��5"��FQaNy�}F���o�9�☕�R�[j�6<��e���1BR��9j���+�|}�j�1I�"�P�����046�["�u��ؕ�Tެ܃/���!*�Ă�ų������[�v�B�������pD�+y�@��5(�%��,�;��HqTA��5H�R�	m0Om&F��Q\���$�#���ƯP�m��������U<�Zʀ\0�س� ������ʶ C!z���}Ѿ���Q�к�f���kulm�3�u�B�y����{��J�D
���h�C52����$#P��!=��?~�/4;����5B������ɥ��y:����$�pg�ܩNnW��4/M|-���"$�Yo���r2ppb��[�H�"n�a�M�%-ٽ74po��H��$br��V��-(�.�cSq�v��.)�G�Ȳ`T//��`�Yk_[a�E��}nu+/��ɚVt�0���%y|ԧx\�i'@�ca^+-�++(\@$��Z#~G�r
���LmQ�8C#�<7� �M�OHn��Hs��:kk������]����Է��|QTLd��{U;�"�]opo4��9g�J`s�a�G��@�V8�K�j6p�o��:���-�K����x�W�Q������K���_��h��Mó��u$����OO�6�@s��d��/��yVA[�(h��fFAsp�z#��M^�sz+3�������������}]j??2,dA�c��y=����eg�&���ʷ���6Ć���Q���A%�pay�R�Y�pEP
z����ed��Q��K%*�|��x4��!�G@:*>~�B8	!�㾱pC�@��^0�^_Ƿ�//q���e�{�ek��� ��1l�g�	��=z���d�T�8�k�E�zƱ��}޵ڸ�����eZ��ͮI�g��r��>aA6z۱G�9�1�S�eH��D)���o']�ք�*�����e.�ڋ���|J�)(�dz�WL&�Z{�
��r��r߹?�-��\�8�bKu�0i��&MB��ͪ��^���ˤ�X�����iB%�V��0�Z��L-ƹq�u�8M�8��8:��~�ͭOܹr���=E)!�e��W�v<V"���i�g�N��	�����{G��\�NE3Rp,���Ņ�J�oٜ~nU����$/j�!G!�p�2�K�*�}��Z�{�.w:<z%e>,ȉ�(ec!t�<�I��,�Srhul������V%�TF�!�0ϛaA�w�h?&�yY���9d]ds7lE�˸Θ};�:'��x����LN��xj��%�C��|06�	��z����F��a}z�Y�����^/�"ԙq���-
�)E�v����.̆""�8�ɝ�!��d�\@�K8EFM>�xD߄	���QS�"���׵+��qۈ���
�J�;À�j%���o��I���e���9M��^o���+_w�LK׮,6�4�)�b} �7릎;�?� �G��Y�v��m�SN��J�`l��'!�����k���/p�c-)�S�n�GAB4��̏�.[�bQ3�_�*���a*�䆧���}w��;�q��+u?'�7J�N����oT};����{]�wWi�C�8*�˘Q���H��x���җ���jf�쬯h���^�|>!,�hr���P:]84Ѝ�,+�K^"��(����Ԍ��D����-�^S��)�(�t�`_�ى��o�Y9�eҿ��k��U%#4�d���˃�A)�^Xy�D���^���G׽}Չ���J��I'�Z��ʚ,��@� �	��,�g�sg�0��_-򺀍+�v	�3�`Ø�V��$ݔKFj�L�d��$�5���K�章5oY��;�g�e�ޫRq5�=��)��b�N�+C�)�+a'0&���H󩋊W\�v���a�~*һ���Se5���|�-�U� F5�9�u�E�����m���F#���1VE�}��_iVV\>�����r�/�*|���藄.��W�Ұ��A�}��@�0�QLr��/�Y�]��Xw�'Sm����l)a�.�]���y�hc���0���y�{�K#�,a��<�|��߯XIpD�dCЃ_�d�_w�g�l�V��&��8��Jxa�� [8����F�1O��Hh㉠Y�I�D*���f�/���a�\�b�т��m\���^[�9|[�v�(鉧�/d�R�V�t�`C���6_��v�=¥H�6?m=NWR[��j�ݷ�^�=#Y`�3ua?��v0���F�	�@����_�Q5t�Ӡ*X��{8*
#؆Y��M�{�|����v���KP_<�^ڧ��9o�l�6��7q��|v��d ������D�X5=
�\����ް|�Aԗ��Gf&hxM�˙=+�k�7"F�v&��dy�.����������a�5;���Τ/�l��7Zq|U�CH�9&=c�}��g��S�&�釟�9�G"ʾ'���Įi�[)&;z�y�KT��*!�4�
C5Dr ��$aj!���g��{��
!�}���Q��=��Kt�+����#�a;�
q�P�V5������t���$^������$Ů��=�Z���b��O?�I3ߨ%�]��P8��|��uO$Q��yd����ei�կ�@�ؒ�a���3@h��dT9j]Z�eRۆ�.���;n <f�H5hP���+�=W���F�Dq"ex	��a}L�̙ec��v/�M��z�"���82�6O�����������L�w�t�]���?1υph�[:M� ��~Z¾.R����O��q�dG�<�w��q�W��O�r'j{����J{^*��K�|�J77Ǝ3�o�ޜ��CYˌ�ZH2voS��i73��%\����?qC
~���R�P�h�E;�A�:�Awn�Vk�%�ߞ ���m��G"A�%�q]~�B�s9�آG|��*�H
� t~�Ƀ�n�l��~�`� ։���h�	�7�Q�7��Иo8[_u?B�-N�}z'���Ru�r~��!̠�N{�("r�P~���h)mdڿ.teĽ�k4Z" ��'=ߍ���;��g# ����Ć�JBk/i��q~� 22aP8���H����a&x?z������cd�q���Q*�C�����.Qc:Q³ܡ�+R�p�f�f�$g�H�'�X�2Е&$��MV_�R��6�(l��m�d�6|��Z��1�i�	�[ù]x�Ě!:��L��+�~%_\d��s%؀�)���%@T˘`U��g��iO� L�_u��l�o�v p���Œκ
��@ӷP_&g�I�CXO{��hz55�D�I9?V�!�S�'E謇���(�%����*��^���Ȧ�s~��R1�a�>�M,�\X�q�nH��r�E���1*{5.p�b�費�����0�\�y!�
�(�U���A�Zw��� ����﷝�|k�Wg�@�����ʌ���/V��P���|2o�1oj��v�j��g���Y�����Ǒ��	��`8���q�E\���$��rL�	>N��Q2���;�;�.�C�������`�»"4�Eb�%Jr���Q�5�o��\�=�cr����������QQ�����Si���n�-z���0h/l����;���[ѿ� FXfGj�,q[x=2���IyQ���Z��ȭ���@}\���6����������G2i��[��u�ޠ(�mT��!�:��l>��[VaiF�&`�:bl�I��ɫ��La7�@`$l�bGtxt�0��V2�ٴ��74L8�h�Vg+�q�^0�_/�!n�)J�}PN��uU��Fsn��a�W�7�9�O� �E����� ~x7G�6�kU��[R8뭣��qy��@BȞ��\? %D�ޜ�5��֪��n�y�R����<���E��C��u~; �[F�Z.d�m��@Q����-����Gz�b9BE/��[�BY�lf�؟�|p�k�u�t�h�����b�������y��w9&$�<Q4�M��GUJv�$�@> LI��f��[&��wy��6�4�������%Kv ��[yO��L�0�eAw����UHǋ�Zp�"�r��I����O��R� nό��(�K�m�2�.e��,۸-0�B��ŝ����P�/�EXY!��:.C��n�.�!��R�� �CR�V�
�7А��QP�s�g�'1짨)ٴTd�Ȏh��gt�(�Z}=�l���g�*l�8�>Ė��8�kB��ӟ
{1eNњ�]��ɍ��qf��P������';���)/�g�����M�fZ��_v\3,�q.Jsa��@E�N�K�br���X�5$�kYJeln��P��8��[����Vu9�*��~�%�'�Ϧ)�V��
���I���h�6��
���R^}�ѝY_�iX�;��%�N� E� ���q<W�ހ�6s.i�a��&R��<?�2.��or�U�i����IFS�w'Zۜ^��N�G�,�L�=��S�W����Vh��S�!����o����$"�_9��˪�r��ր���,'��y�c��\!2�&-U�{o2K�7p�.ˀ�6�f>N��^��?Q�Ԉqi��м��C!�/K�/Z !.���)��6�����Cm?jY}�t��T��yeP���p�O�'?D�<�8��TE�O��A(�ڭ��4�l��=�K�>�o�?�7��u7�6�v�b�B���l!<�"1T �<s�ewE��L(����sJ&��wW�s�J߄V�Z>�ʒ�f>>5��pq8|Ӯʭ�p�fL��l�8n���.�]wr�D��L��n�`�`q�E$����v���yd��K�(�[aɌ���ŉy0���J���+@�L,�T�^}��Q}Q�����s�EG�H�)��RJ�`ܑ����nA���!�H��pUå� ��;Ǽ�Xl���&���$�̑�	W��R�s�E�U6jC�f=�v{����K7��/����� ���k�x�̒�T������%o]�pF��G'w�����j�D�H�Y���/�ï�u���{.��!��-'�d�uBQP���m����X������:E�I5`����W�#HxIj�c'	����A�G�K%��}"�ħχ4��_���`k�j�Zv�C�w����֬:�U�ᑦq�x<�8��~�[`��#0@`MwbЗڅ���-�嶐TkR`WuVj	�j�b��(��&j7S��+�������y�q�S��<7�G��rW\_y�`�����o��Ǖ����o<�>Vc�1�Cy3�>��_[���bFN�DG܁}�X�}��\)G��t��n�L2�؝&��c�;�4�Kf����Xg��h)�2������X���Ό�0nMZ7F<'6e�����5�h�JKf
<Al�����/T������1�;x�S�;)����s�^��oH���[2m{��|���,��/��V��x�3�;ĭΑ��O �������݉o��Z�"c>`Q�"������S��<�G�3�j?����!vLZ���?���-= 4�ۅ�a��O�[��$͸&���U�Z���� T�����h\�^�	G�Pgو��9U�&���e�h��Ow�6&q1�R/��Z�-pK�h��ǎ�ph�St��$�&t��������h�_i�" ��Ha��.ü>f���9�;OoUT����wڊ�AN��I�������h�d��N�~�zM���� F�q���f�RH~p�?�6i������!�����ю
��nJe�X���_��֞��:؏,	�po��o�z���D�{O��c=%M^�T���\�t���v�5���+;_It�#�
����쐪ݫ���V{[ɭ���m����3�m��P�a<�"���E(�;���@��"
tH��v,>Ȼ�+�Őa��߬�%̖w3��G�]��B��`�t����a[��W)sT齿4z�}���q�����%�*Y�&!a8��� �c���8nCBG��qi��X�WG��DY���2g^�8��j��hи�V8ѭ��� U�;:
7��.�Z�U�fS�Q���nFn�ll��<5���^1c���h���2H�!"wi��tR��0�D��b��@����0��ׂH����^�����/����S̶{��p넼�YE 6�c�쌚7��o��V��	gL�
q�ŉ��iPn���;r%:��v�a�s�~�b#��C(���f��ӛ��@"�x����!h�0����"C�q��L R�!,��O�^�yE�&F���� 3ݰ�y![`V�����k#�Ħ�2ց\�;�
f�9m���]��S��%��̲܂+.���ϕ7>�Wq }~��fQ�n��Kɞ��ɽ\��p)��4����ݛ�!N?w�K���G�M[�x�`a<���%�y�#��&�>������b��Hp\^���)������C�����N��d�l�bL��=OM{xvћx��K@Kl\YH�x�Y�!Lg?a����� �|0:̙M�u�4p�"<g��:<#p�bdl���ZR��`��b��R��.��>�V:�����Q�+���U|�Ak����>�C�L�.�WK��lI�j޺K�}�����p+����]���=�0=.0"%\����#�''�QQj���
^UXF՗�S���P�Z 
���+�v�д���j�Yx��N�F]��4�H��dO�|���w�$ʒw7�:߉b�g�Ê�v���cۆM~�̿JU螳V.�^����}}��`V�Ø��w�[��\�rp#i�h��%\����=���GqO�ln�Q��
�#TlfxD���8X��q@�8�%���_%�2��?E�'�����S��m��py�
1�������UXǄٵ���? ��pf7=�R�
�ZuZ!��c�Ȧo>M�W�u����N�3K�E�*�v��g[yf��M���j�&�M�^�u��/�L�2��M����n�<ǪKZ��D���M��$O��oI$.�^.����5��b����8�.���ׅ8��^݆27/܍����X������T%Trû�
����JF$�i�1tZ���C� e�ܐ�5� ��5VŬ}��&瓃v�N�9r�Y;�Z����c�ί�lj8��Z=��<��Iᝰ�ؓQFL�}��a�S�N!_[���[���ۮ `lBH W�T�f��|bk�$�"fj��Y.,���-�X~���X�yG�k߈��
2_�P�h
�5�8����'3Ǌ_:�s�x�>/�t�P���r{5����u���'5���-s�儵�<����P��]<A� ���r$%B@�#xH�RS��N���L�r��}�7�X/�����M��SpΐR�*�=4g]n��q^��٦���\���w���n��U�F��tn%���E��>���V�&�lۨ�߲|�M��[�!X-f��q��R�z�;�Q���l*ɞ����"��PE�ڗZu�����|�G���/�G�D�d�8�k��9������s�\�#�@��J����Hz�y�0�cd�ʫ���Y��C0�H�]����c�t�&ϭ��EՋ?���:tR�?�!�w�&�vN�>Ţ׸qc-����FA!���.�wr���Dd���Ӥ<��� 	��Ӊ�+	�X0�P�s��5��l���$�N�iFR��CU�R��k�<MƩT�6/as�~z��4��6!3���h��N�k@�Զ�y>ۨ����u�-�.n2��c�+��eQ�䳡�%֏p��F�bw���ĳ׷VX	�,$&�CP�����m���I�=D7u�Z���k(}/��G&w����~�4V2�d$��h��7a�<�������z1O��t�4a�F�G
����uH�.�I}N��6z `����I���z���u�5{}�4�c�����C�`�ƻ.�!�fOq �{�9�ً�6G�`��5�JǢ�bs$��թd��<�f�!\���,#2�]�.��h�OP���鐳8؊�[q��w
8L�n"�0;6*P�V��Z���q�L%�!��{B�L���^,]k�(B� 
���I��V��e��K�v�Ȧ(�!�ӭ8�Y���j���J��wsT�$Ƙ���L1_��;-mo�s��E)o��g?�U�9��3���6s�rU�""�\No'j&u�Kx\�#�������9㭰p��e�����2�έ�96q�y�O�YK�[#|�Խ'MF��mh۞��'<�@è�6e?���E۽y�{�ā�2�k: �0�U����Կ���T�Y���8D��0�Ĳ�`��
Y/�1ٲ��m����К�-[6�v��twG�$D�V���n�N=��/�N�v��lp����l��T����]C�b[e2���g���?DZ���Q��r��SěP���h;MCcX�.����Q�C*������*����?Ӎ�S=�����(���h()|-�x���	F^h����]
��8��]�B�B�7N�<��o�c(7O#=3}[�8Z�b�iX̆V���4�'�f�/��¢]T�s!�)��0�[_|�%5��.�ݡ��,�βF3�8���%��#�P��h���i^ٶ�}���q��K�.�t��c|~Ck���g���/A7��	h({�
���ߦ��Lҭ"8�d�9��2k8��H�vR�%�e�w�@K�W����Rݐ��|����əX��<��6X��
0�z�$�?�T��~Iv�h�t��N���Q�%��x됏��1I�kK���L������nO=ë4�z�j\��;,�_��&T�� u��~S?SM�Gʹ��]�&ՠ��FS���8��`#�!��K���V	�1�M�U毘;Ÿ����@���.�4��oXU'�f.�]7�Y��1~:��%*/��E���%����7�K���Q/�摯�BW�M١~S���vKLvԴ�:��]Y���)۠Dj6����)ш9���-���������I �4jj��Q\�Z���k�Y��3v�|!���U)(���3�L�E����F}0&k�p��0B�+��o���g�qC
l�����q��c��s���^C�&V������U�K��7Ε!���$4����1/����#��0���&U��#�7VB�����c��,S��Y�^ET=ĕ���roQ��e�4�ڐS���.en�'*H2�S� E=-��Iz��mh	�-�#�FK���$�U���=���T` v�h�ɲ���OT.(�"����1b�4��k��/E�6C�h�6�xQ\��쫇��\u����mŔN�lР����[���ɹC�'�(�@ڇ�����������R�9qY]���h߰r12�P��Æ��0�)o� '�s[��	�V��o�%�B.���Ze�\�f`��5$?��'N���t��%:�5��'�����2����ܱO�	\U ����I^?�k�������D0�Qo:#ATF�_$�h�Z<�{%_}�`NA�O(S�2�lo��ٯ~�8=�\��Vݬ��,�v�D<[=t��J8M	��%�t������Ϭ����B!M)u)֣D�P�c2g4�M0��
��Ȕ������v�%c�
A!����bU�T����Df�*��p�A9(<j�.� ����AG&�,�6T !�ن�tV��;s�Ԗ�/��xI��BzT�3YD�4�!� ��h�d2א���bLX��軬ٗ�)"�3+�z�O\�ɪ��L�u�l^D�+�)iDF�0��}+3��PO2�k��(K��WU�������A(�2e<@�������t�ق�T&��U�y$�16ȼ_�,�������8z(�2��/���?2���cT �I�N �:s��`�Ƚ�P4�-��pa��?��6���;���0k�M;nw6Jo�<������H��yc�!Yʹ���E]�x��w��7>r�(��AT��$c�#W���v�J��X����4�ps�?��Cp}�Wd�ȺW%;��9q1�װ���'��	