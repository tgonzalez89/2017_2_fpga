��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR���[{�T���CK��TC,���:�
&��d!��]9�'D`�"9 S%�aQ�`!�6������V�W�l�a锦E(�\gC�slu�4U5=1�N�m��l�9ў��P���B�@+yg��=�}|�6�`hD���PwҾ��h����;'��P��,�cZ��w�+a���N�sҕ鹻qt&	�Ny�>ʢSi�n���;x�T#ݿ���t��dQ���C�;7��!kg@D�=]a���2�Li|�?_J�]�L���ӵ��L���4͓�y5�k����d�[�K�
M���H��U����p
G���0�v����-��y���|���,�E�G��	���9��s3�{rS��5bu�3x�	�_B�1���5���'������;:#D�31xEI�[�q1�':�- ��<AB=�Ii�A��s�������`=H� ��������'��_QS�� ͅ�HP�u�r1>NN�ӆ��wյ��KbcEǉ�3�����'JqA�"nſ�u`��9�O�>���'�����UZ�
����j�ܥpO��n:�६�X��-����W��nX��C)%4��o����3*�j�0�)�q����{�`����Nx�Tm��7��o��|�V��T��a^Y� �����>(���ǈ�)|}�����&0۟��x�)+��}���X-ҙ�Ix:�sM�5#Vq�4��P�L�W����h~D�wP�,�^�Y0p�b�¼uoͨ���K�7;�`ѫD�8������<����H4n�%hi^��m�Mp��rr0����T��D:��1�3�ަe�Uї���"�J�x	���S<��fR���?q[�[�L�)�����X=�a,��eTd-wr�lVk��#:�M��o��:� ���iNN��Z��r�\@}�������[A ��֒�	��k�!���N�9�
LL���;�8��\�W� 0�]���0�(��7��a2�m1�D���'����ڇ�U5���]�D5/ˈ˰�b�*��.���$� ���d�K~f���[Z�\ߝ�#�]:E�B�ur��H�,��h+��whֽ��xQv��F�X�#Ѫ�v�٘Ak��خ1g��	6ZSV4A�(�	$c�GA�9�ʷ�^O`�Ω�I:Z���D���P���ґ&��3���܀��0��yh��Y��2bWe�Vb��9���5�#�0AբD<���2���W^�U<7O�p��F!��u�a�qt#0`2�+���:�f�Hx�j�a�������U�w�➏�u7Q��;Fxp��db��@*]z��4�C�p���^��8�!���x<��D��;J��L�ˮ�J�
B�ɬ��\^2���������v��p���v��my3g���5Ht��C�%���vب�.�E���YLiY@�񅿠Rf=f�ڎ:+ ��1Z��@�'�-.���L�8*�@eWȓF��1�C�鹦O�y�b�`#�j�1�_�GӼ�*�y^�ʃ��Twf2L�?�F�3��!�@[A,�$���)p�w]���*�a@�g����n|�������ѓ�p�mU�E�֔j�/΢"ϋPx�d�M�I�X*�h��a㚊%�jM�@NTh�u���"<dY���N	u<�NO��^��cB�ߩ�E�K�'�mo:�&c�g��k��E6���Ϊ�W�ُDMK�w��"�Ob=�juM��;eȥ���B���9��怅gٯ�G���QՂf��I�����qV���z8
�8�ޥ���w�&��j㞌����qEOoï���'oqT�_�b�(��mǷ3����	�THιB}��C����apz�3�9NRp�\�2��C��kl�"��texୀ5���*_�H-HJ�kx�ڂc �e}�'�\���(�!{��x,����Ȓ���>���muOQ��r�����/'c+@����_ہ�3�`/9�ɂ�F8-D����pyry��DWF�hk�iz%���O�f+~�έz�p B�����J~bS�G�h��3@�0��AF�BA�� ǿ,��b$�W�����y.�B�T��	k+ܮ�?�߄�wL+Xl�*R+��u�U9t��o��A�E���H�hB���!�M�)��{lN$�B�!z�s���˾�byK} ����Pwn���D�W��oc_J.���@$��><�؍\M���C̤�}���);�3�X-κ�@Ї�7xrp+M:k���@NU� �lw�D|�r��X�З;FM
*7Ldj��((��7��+������h��=��������)��)�1d=ɢ�)��yW!����2���J .@,�mι'&��d���9�D��o����~c���`��M�0��y~��Ӑ�����q��}oq8�,��׫��3�ȤM�ދ,�?Iژh(^M_��b���iD�&�Uk��=f�CT�:M��4��@h\�JNT&�q�.�tW�%��"���q,��_�!$�N-���V��e�?�Cu�R��J���z" ����8a��S�x(��Q�E�]Gt!��:���Y֘��|r�K�8U�(M�&��GU�>y�?��@�o���E�a ����GD̗,<Qn�,�� wu���ȋ��m$����
[O�b��%1�_w����S�Vo>�J��)�X+��T�J�N �ȟ�	s�_�$	�+�u�Í�x�,t�|^
�O��h��{r`$n~�5:��oa�ɜ�&fVW�_ݕbۛ���u!��@�X�̴�(�]�ڡ9i�/�*k�xZ�M��*_���D�Bd$WB^��dt���'[���y���,�A�~R�E�6.�86��w-ρ?{:r+gj��wI!3�8��ro�G��
�q|P�G:9�C�%}"Υzh��Ԣ�@��{�P�z�o���"��pfkl�k�� #e�;A�z��Xlg��K$���{����{̷�c��G���g8Z���(?+]�����*2�P1ҥ�Eiu�g���J��%`Be�n,jZt�*#H�/�ַrO�0A������ӳ�3w�]̦���f+��FBM:�cƂY�P�ݓ8�����%���}7����!������C�e��fRA�	U�Q9������Cq��]���{�d�,/P�H[Dȫ�V�cN��?j��@av憏AIHM�&k)��!�EUA��Qk���u�Z���\q�L���ϭy�B:K/�:����[c3�Sp�����Rz���wy;hgV�J�e�J��哒a�������L����	���d��V UbVY7�KQ�H��*�ox	"�ۺ���$:$R
�����!	�$��W���3��:��N�=���{y���o�$&���~�k�E��51NȈ��_TwE�V�ڹv���������!��=�q� �t94����Ľ�b�g��~���f�v�����sp����}7��P�(W��p�f�au�H!ߔqM_%B���U~m� ع��k3u+|�Y�W�FB���f�H�\vJ��HB���ɸ�0����l�m��̌��5�W���!	Dz�j�S���m�+T}�P#�)�M�������&*��觻e�@A���J��h�K�8���X�r7  *�ޛ�IUyQ�۴��4h�=7z�Y�Dn12�A({pr�2�cv�t���&z�g'~+0���Ő���fz5;�a7]zk�̄�ճ�e�6�*P�Y?��Oˌ��##2��QT�u��#��/�T����Z�{�k���t�x�w �ه�	D'p�;��Ld.�T�)��h��z��+ӋDk�ΐzf���͸ts�m�?�Ş�x<��e��/ƟL_f�GD����`?_~/=U�����a�)�yf����>c�����2��N�7�*1|B
)6�����%k�8���$�9��Dª��[?W��s3e-qq�0 yv �ާ酩x%�u�-g⨻�V�1rn�r� 2i�V@���v;�ɾxG�4���h���T�|!G��	v�	�y:�6�єV	�<M���;rk������T/��#��L��L�0����c�v�Y��MD��Y�IM�2Aài�����O�v!x����X�z�i�^��Z��i�ja�(�I��=�ºGǭZ4(7�+��4U��p.��l��ȲE_�m�͙`mJ
0� 2'�['��O�#\��;Y���*Ffs��>
�G��¾�!xnA�y��G�Z����~'�7H���8i���V��
����h���pzwׂu���QJ9r�qfZ�u0m��v�!�s���6�-P�֟�'�^���3��O�>Q��"G����~�^I�
Sv�{���u��g	�f�\�L��.��1����a�\L����¦�2�g��?�3����#�����d��Z�	Z��f�i��N:0�;��������3tHS3"��>�<n>���`	?��z����+]�v2�knOe8G"��#bq�~=l���Ng��ͣvS&��J��'R�gL	6p�3g��<�{�\�q��Ew�S�]����h�?[�U�ҏP7R���A;&r��0o'��Qt[�Y m�·-�����^�o
b�>,m�p^ ��M���6���
2;�|���Q_:e-�[�Cg)R��O�L�}�h��y'm6� @�^�N��`|,n}5*�x:�l鴘䀮�0f�4xe2�>�S�(���)������m��\�'|��Є�#��^i �V�:��D*���62K�D�k����§�-4a�U�ס���&!MyT�5�{��8�!m��9�@9λhv���,��]������VV�R�f�k�ě<X*���� O"d2~��E�u&*�	-��!�������U�(xF��4WrY�V�E��`� @>��p-.4̣DՏ�ș��gV)�*9��d�#Qǌm�	E�!�&�ѵ�)��b��e� ����H�D��eGR�E�s�T���pA��X�x�'�L$c����&�����Xc�-�%�H( �qP,�w��[m؁�hz�Ӗ����"�1����kNVM���va�~_L�耫���̸��k�i|�5�X�#	8���|k2��ahi�z�J�V��8 %�����K��D�1�v3hPl�p031�>��}���Z�����ˡ ����+ɞ*i�)��8H�܃ˁ���;P9��֖b��ϳ�)�2�xK�_:�۸�z2�j�;j��Wh�@$@��褉�l-;�f��.:��>��jyQ�*�6s��`_ݳ�Z�}���@��6~���T�r�K���9/o9��P�a
��2��XМ��
��t�p�<L��.T�"�s#��d�� C��������t*Z24 �F�c`��R�Z�|}·���=�����p�P$��Z۠}�9AM�@��~�y�����F��:���6KK��#i����Y�L�Mт8<;�֎=6�t~��X�G��^Ԗ�"�)	��\z���j3�xIҋ����!)�η�������k��-�=�Vy9)�H�7J�[`���̼㽐�3��V��&��5��Z'/b��N��>��=X`��J���1_`�ݐ�:��0E���lV�M�b	�-��Er���q"��d�0����KH:�fS������ȶ� Y�����d�T��Z��%�d��P�)r��v����m6�D�f��5x�:������L4��u���Μ�~�C�7��5"�聆-?ZO��
Zo��iu+`Қ������c@F�Ltc.y�]њ��w(���'g:ȟ��J�9�n5'�l�G��T��ӏa��k��<�m�Jb9���J����0�����oao<� �S.�b���K-�,!zGU3�J!�dT�X �����;�3��!|D+�g�� �cU�c8�B���sf�$E���X�p%���-+�����]Xq4��A	�Ŏ�YJ�lU����o��^.}��+̰�toMd򭀉�h���G����4�����(G�|��PU=�����ę�zF}��Cd��<9)M4�����.k����ot
�+��h��HF�4o=F����������v�/;#t�r�C(s�ۋ8�?-�Û�o����q	*/�B�c��q]���Ŵl���<-�1�yl]�)N�����Gᅥ��a���4x�,˃=~\ܴ4��!��1��㫆t�������z'>0:�`��h+m���H��۹�a��Cg�.�����۫-�o��Z���=}" �����x�e%'�Y�0ٶ^7�c�Z�)��{J����u�v�q�'VV&f]8
{�O2��T|3>�k	��c�*� Z��a͟��N�sV��~N��x�4��s�K�d6y�CcU�ܢ(G.Y����f�&P71�q���T�����h'�:PR.D���4|�UA�'f1yR7��!c�|&?g`�����W���SO�_�|��0�*�C�b<e���s
�t���߱8�[��|l��mK>���F�"�->��њ��.��t�x�9~6ހ{�N�e@�+�(�'�����hC����΋ @����Q�&&B���b�_��8Fw�j]�[IY�(�E�4�;�)1�2��#�'3�iy	��hHB�G�L��S�lC��.ykS)�-�In�&奫��h�Z�/� TcX��EI��"�cW$����P|?ᨋFO�[:p����.��nTIR=�x�ȝOjU�'��m.Y�*G�':���u�ܞ�!��$%�@l���<a/i�W�y1XE���u;4uy�p=��ś�陣E�!�� Ȗo�{�9����̼z��(Nli�%�'|�%g�N�׾��^;�,�"@�:ڸ��{c<6(��a�N�-,]����x�)�� ����4�����'iʭ�bp؂�����MU�?�G�f��Ʋ��LeA��Q
fFU���G.��'T�w����j^�lja4���=:o�efi�y\@X@�p��R[�m�f����nܦ�zLh�g;-�T��{�I�V��-/-�#X��{m�-߭w:���ֆ�r���ww����r��Q�Y*b��d9����6b�z��'��,�/8^����
��b4��9	�ݡn8.�S�y��J/��j��/��t󲿙:+2T�e�:�����ȰFSf�R	C��"k*	pWw��q߀����
G��f"(e�<�I�F[�'���c^~L2|�as���o/�<��cos��qf�_�?���2�AK�j�)�R}��̹�B�=R����#���O��<�����ؓ����Р}Q_=?�6	��q*�Jc�(��
Ù�}�?���K��!�o��y��3��Meu`�1�O��C�6��Q<��V+z��ϥ���T��=��>~V�9��R�i)E�xm�Aa���ZC��]w�K��kFK.!�	%���\y�o�>B�35�I=����0�������
/��H��Џ����M������
?�% ]���U-LZ�F���r����U��L�;PM�pu������?�� 