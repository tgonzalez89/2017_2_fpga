��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR���[{�T���CK��TC,���:�
&��d!��]9�'D`�"9 S%�aQ�`!�6������V�W�l�a锦E(�\gC�slu�4U5=1�N�m��l�9ў��P���B�@+yg��=�}|֦���ָJ˰�E)!5���I���r�f�IT�A� :�����m �9��0b�Hi��e�P<C������v'�^i3�(���i�(W�I&{j����\�m�5Jl|��Z&��g<P��������5w40��OZ���򅭽�㫷��"�שǚ`�:��j͚0M��w��()�z4:�-�V��Fe9����&{�x"p��nQQ��kn�;�,9�ڧ�%�'����ǅ��^[��F�8�!,��MR	�ɣ��c�T���zA����D��R�;�(�۲D0�I�2s�=Hc7�Wd�/R���!�������7Q�6j���d�&l\�|v�_*:��M�O����2��A���z'_z�3�A��z�9�$4>���)T�Xm�ۡ-�e�� �%2�# ��1����Y�D_�L���m��ɿK��RwSn���¥��RD��)�Y����0u"ԯ���g�p
L�î+�����g�6��c��*\ù�D4�O���Ft`x�E��Y0�0����A��b(Cx�]2h�9�z�@!�y+��������^MQn����;��4r�p���[5h5|�*Z��}��H�6j��A��w$/s�[4qG���f<��?�&�oZ�Ao~�X�1?|W6�rŧ��F����Ѧă��V:v̲⹀
���������X�D�$�3yi���N��e�����al����rrw�ҠS����Fw&p�__Č4KW� -9�N��>���y��L�_��hW^%�{ҹ~L��,�D	�2*a��� T'p}$�ǯ{��֞l�2�<���o�޴9�jj�u-�]"��L�l���us��5��8�C27����Dg8��k����a���+�:�P	w�'�n�̺ƪ�ߨ�hJx�E����~�q5�t�_�g��W�P���5���Bk��:K!���+�8�{-��t����ы��§�#g��(e��s�V'y)�;F>��9����zێd�x�_J|����r:Y;_��E��M���]�� �blw(u�����h��AS}I,%`���ǆ����Ϡ$�M �Qs(��u��Ǘt��A��E�*��eI�ٚM�e*M�I�9��E������s(8j���QA����z�D�'=��$ lUV9�V� ��@�~��ksF5QN��c����JZM|&��v�H���C���@8d�I��h��K��V��wi@��>�~��P�������y��#��|�s)C���M��mw���l��B����C��^ǣf�GE̖`�~��}�@v3���wv�U܃�����!���C��G
����8���{�B��H�����O����p�&�LƆ����42�\O d�'����!~��� dF��bEc=�J���|��w�%�A@��J���ob����-^�r�b<Y��e�H��4��-�"�V!jO�Jw��o�$��{W�,(i���Ʊ&9�ҟ�����@�6���ys�|�{b�2Q�!�v�(�^r��Tb	#�h�b��p�γ��)���R`$`�!+s�l�b�0(�{�ذ��rs3B�dŰ0n�`O� 樼���ˣ�נ���a�=�:-P^�+J�w;�yC�:���7�qv
���1$�ѡ�֌�}�=�[t��W�c��
��S�����0S��3)W~��;��P�`�4F2=��¹���17���0�V+��}T���ұX�����T�Il��\~F	�X��e����ȿ�Yhx_VQ�r���V����q���[�O�p�Q����L��A�Lo2i�����c�3�Qhb��yze�������I[Y��n�����*E���tNV���❇��[����-z�-��ol��ʹ�z+2GUo�~t���$���]42Q\G�!����5�##�RŢx��z���!�1Fo��.��p��0��A�dbJE�>y��]_�v���"��;��, :f��a��E{Q��=���к3�J��$6r6�MƐ>��+g4�T~�Ŋ���~���n�Ө4)�����Q�����؆L������[�a�c�ү���h��O(5�2����[R��"J�"�oޡi�(���<�ؕ$��}��ٖ9�Pb���XpM�4@�	���;��rp׏c��IcڸOy/����۟kʒ�@3x���V�:��:���@û
;ʿS�|����v;�.�������y��X�1�k]�`�+k�ö�=|�[�H�P0�[2tL�T������1�NwSv}�S'A����O�s��;�~w{]w_���$}nyw��puRq꒼�)�tz�?�_g
��KE]Y��e?���ӎ�Ӓ@���L��ZB<R�D|��_�?�C����n0��[@X3���P/����KO_Y��T��|lܘ�e�D��)G���rA�z�s^��v5��~�����o��ݏ¹R�ЭR�,�fq+������[�T��J�w�Ѵ�Nt�H��`%��j�ܿG��
B5�W�D��js��R8�K{<%A���cuk��p0pw+ !r�A���6�cU;���t�y��B���?9��/��~����#dSJ�������\?aD$�"��Ԁ<g,�F>}�ډO���ܮs;�`�m�
#mf���j��/�͍_�b���`�om����q-A���P�(ye3�Â��ZWd�.��a\qf4�)�G���c��B/P]���d��=��^m��Ď�4��J��XX�S�؏t9*�+/�� ִ2�r���:����l�����t~$�Q��L{ǖM/x�6ϧ��ZS�}�����-��SN�Sr�>�16�[3=g�|��z��}fB�4��̯k��F�1��:����$J�&ɤm�O�����p�������C&�Nj#��l��XeJZ�@
!!�$7w�P�G����S{ʲ!}c.[^zdС[Uд����,/U�+ �!��|zq3�����O�^����ːG��d�P�>���E���o�	X�[����oK���Mg䵷���f��^y�#���,{ Zt�rOD��&�"�j2�(<%s��k�q��o{���9U6 ���|������vC]j>b�R��kcӪ��ld/Z��D x����f�H�}�	ō#7p~�Y�������/��nX����{Z��6���k)|�a5irV�C�:;��`:{}�֔1�Q��� ����W��dL!�t ����C���W�pg"��`%(֣"�z�?�_ͷ*�'��D�/D ���f=<�<�zY���u;p�r�MS�W�����̳��^����`���i��$T�(2+G��7\�dB(�V��,bZ�8��L�z�k:�xC!�ZJ�55ߌ~]e[w�=H��P�w�r�nU��P��I#:�K���0׹�*js/΁�Ʒ���8\��Xۜ�
�_2cTB�ҙ�d��U�n�p�u��&��N䘺�6��#�#
���{�G5l`�	��}�7�1���U~�\�W �O�iZp���� 7wJߓ���R���N9�oY�=��l���t����ۣ�-Ǥ�W��D�<&�(HZ��D<�����ڷ
�� ��CѦ���ș0%͸||�U�Ð,�dU��Π���E�Df��Jޣ/T����+/1aiO݊��"�0���wۭB����-N�|�f�6�>"�k��T��_�����>����kX`�Jw���ǻ_3�՛{�����4�9>ޔ��tO�(�J�f&F�WJ��m�� ��+�o�5�8��+`��p!Z7�Pw��mre@W�!��C`pjX�`����������A�ȿ$0�'�Ϲs�h)�&|����/
�Ŀ$��G1��6.r9j58�<r��t���/D��ЫdG����5��/�q�Ss�rE �7��go`����Z;��<�봊n���ǃz~�%�B�Ҙ���Cv:�uw�����emLf��d���^��L�}�R�?P!9��w���N h<�	pa�h���m:�mKqn�b%ǿ���
�(�QA��oG�'��1����h�҄�8��,��Lx�G[)8e;�?3�S�3Qa{�#E��Zec�+V�c���~��!�w�<)*Ǭ�Dм��\:N���l6zuښ}g�� q�.��'��d����߳��݂Hz?� |x��w �=�������I��;�v��&e�e N����x_��W��7V{$�$+��47�����Mip����`9h����FZZk�5�<��θ�5��{�8}�f�n�6nx���ʔ//1de����K�;�rs�_�H�V>�\���Rb�-v�ޖ�vy����Dz"�5-Pu�MڱrG=q���l%�	������&���Ϙ�Z�L��`���e$� ���m�l��6-�9C
B���4)
5aѿ��Gϓ˯R��]�ՄX�ӽ��ĉ?�IC�qc�����k%�r��b��t{gU%g�`)V�K��W�R_a^�Jܢ}؊w�;�O�eL��#1�hV nn��Ǣ���|	ߓ%7&�U{�@�e�!��ecQg�v���`��r*���v�6�- L���я_,�.�mv���J��:�hG0���u.��7��](���NW��^��ϡ3�ջ!��2"�ŋ�)�+�=�L�6U#\�5U���{�/����܍qB��� �W��˖��]��)<�o)���t�vW��i��7JuaT
�T�Lo~Y��p���O��hYeO�d�����vB�!*���r�S&��/QKF
�L6��+������-���iQ��y�M�cx��te��}ѶB�����h��� ~�iˀZ����v�6�+r��ng	ۼ=��dco��s��&L1� �[aS�;����~��U\x���Bp�t.�po�H��-�j�dU�KG��	��3~y�Ź_�w0J��\b�kB�w�Exc�e�?\U�be���Zr�����ç,�^6�!_n���Ĝk��23�k�bY�ʟ����,ť��_Fơ芥J#S`��>wD����7ä���1�ܱ�mR�<b���̿ƪ/W73О�i�=W���� 9��w�)�P�Yޅ�U�R�]Z>Wue�}�R���ذ�	��3�f�TCb���v�R�ښ���ۈ�!�����������
��R�@͙�"Q�;��$�������]Ձ򖲿.��+}�	<�\�2�����E��@��`ť���	�/D��i��joo��|	kﵩ;��h�1��ס����J�D�����x�j�:��
����,> �I��sw<℃��#�y���7[
7M8{g-��[sj��a�k:jAu���c��?��a/䏘��T¸��9����L����w�Njַmd-�����mX{�ر !��~�Y3v����{̸ͭ$ǉ���������=�̾��۬K�!N9�g��xš53H+������\�m�~�r��~�T9z��I�885���T(1�#v�L��?�
{�ʨ������oK+*`d�	lG��b�5S��>�	VA���\cl��vv3s����
 ��K?P�[rC��gA7;�O��L.{�Ew\�
k����<6A�_a ��1f ]s�S{w81g���8r��Q�rG��o�����>6zbx����,��F�5���o�Y���jn-U4�ݒ��E��K�B��T�/K;�����뼫�9�  �p�r�X�/�����5&c_�V����6�6:�vm/z�S�fN97�G�gt\�u�����L�wn�͎��"��ద먈.�y�$lB�	`s�G*�&ê�)�ו츍.(����ֆt�q�(�](�F{�+$5�кT�2]i;1��c������Z����9N�j�kı&t$w���?B;?��Do~g����|*JA?Z
�F�["�6�)�9A�ٴG�|�L`��K҆1�T-�d����Oc�L��'*Hf��DY#^�!�\�E�2~�� �ʉ*�Q/ �2�_o��J��$Ϭ'��r�R� ��yV���� >0�WLv?�u?�:%������Y-<�=�����T���_�3�
xK�X5�!]0��
��،5�y�L�$DfZ��=O���&9q�d+���Z�g��ِ1YW�����6 V����U���9M�Fޭ ���D�vԀ0}*���Ej���C�ο�b<�����ycx詬�
�
���,*�ڨ�� DF��_x�rP���Fm�w��9.bR�*��BJ�W=_əj����p������v۸&�:'EkJ+����'e�@�ri$C?z(�w1�qL/�^��n1&,�8|,����3�HKig��x\ 08Z����rĈ2���5	�?�@�_�npȵ��%KNOj�)+��/H��6t2x:E�W�&��1b���� -�	mڌ���&U��k��� {ڝ��1�	h𒙇$�?���u���^�)k8�ZSn?���@cx�D�r�b�4�\˙�<|�W�Q�����
���V�l�Ӈ�g/�#TC���끋�A� �v�}$����3�E� ��g+����T�\��~��KC Z��)Nd`Pڌ�Tk����|9��f�����</w\��~���[�2`R�n�︈�h�� �a�� �ɏ��Dӈ��i���0w%����G�<��?��55B@A��Z�]x�Y�JL� .3p*��U��
��R=��7#���N�|�[+A��s_U�5<�k�H�ֹ�թʿ���J��4�Ԅ���8D%�9��ь:�@	�����D�P��h��G�3)��aKl���r	��������1��z/Բ@�m����#���߫�
6�������D(�պ�x���NVG�E
l��5ԝ3�p��P��z��ܥ�">���ir�Vש�\R�\�.mh�j��`�%M2����n�?����Pڵ��I�)��`���P{I�RE^.]�T��˷}�AM8�^Ёk0����稪c�R* q&V��*��$������	���4;�(6x'��qD��c��
rb�����_y��eWZV�(q+��?��5^�4F;0�β��[�ד��"�/��,_�9��)4��Z!l��C�\�k���k�Tr<ؑ�9	o٭���hG�J��b���оf�*/�	��Y�7�%�K�aI�����]u���[�y�}.If��6�|5�X�m��3+`�
[���dt��vM}!��`���sWe�cȆ�-�;��B|S�#�hɻ��D����d�I�����%�_}y�� ��=#��B��ި�>T
������;�~z�S=\�����a�7J��,g�ģ�D�B�d�r@'��?%3����l	5u�ڬ�l=Q�o�Ѝ����-�k�`���.$�E����w-��:E�s*`�!qܼX���KNW���`�'�Kc���BN:ā����F���������,6�ծe�����B)kZ{�� �.t�@HX�0�3	���GI�"��M��X{��];e������l�!%W��,
����c���2�H�So����䏁��*�ۓ]<�쑟CX0�v�C��ӡR�Y"��K�+Q�#�Yt��K�SC�<4p�M�1/b�~/�ޝ��A����y�Lc�;[��b���W��p)�F��CL-����fy��Xai�*9��uWF��9�T�X�5�ĕ�y\��p�_ýUʒo���>Qh����fuG��?
즥���mgY����
�2�#<�A��&�W���n�)My,T�ɫ�����1�4���ۡ�Y;�`�8c���p~�C���a��g��{����FK�(D�pw�L��]N2�� \ݹ�$�w��c�zΦ����)a��<�
����5_�٥O�6^�Rģ�Y7�7dF���-^I����w%�^���7��ܵ�6�
m,��YN�0<1]Y�ف:�dle)�W����y�L��8�x�̵��	|u�U�E)%G�y��_�Bqݫ7�`����,�-?����m���:63q=�neZ�-Q��c9P�_n�#�J��d-�q�z/^����8.�$*J.�X����,��l���*�`�H��ttdX���sЂa_�~�QF,� ���m�a`�#��������֪#+�C�_H��.R�������t���h�bF����rd���R�������x�T�o��A�,�\�>�]�8l�P������������x�Ε0 I�@��Q%H"��	"��9	�䩥SV��6FY=���1���M��=}H��&�N���/�=����S���N��[�����[��4�F"�Kܛm���M����e�4�]|low��ƨJse�[6���Ҽ�p��O\'b��h ��<�2�[����a���Y]��pi��[mȋcm�ɻ�υy�Z���Pڷ����ѩ�����g�|�R��^G9����rV{�I������M~zFEs��������>��o)A�e��x�~G+\!�g��������H��A�=�N�S�|:8��*n>�e����j��yT!cJ�ܺb�ٹ$���m�7�÷�����f��v����8����0�AaF�%0�3w=T�U���iS��ɹ�b��=��~#�[u��K�����9@���������C2-�f��?m�}�� B��TШ�U5j__�&�%���d�6��8��mRl��?�5H&#�<�zZ��c�"Po��I>uX��'��R�y��r���B+�$�5���pT�����q5#�}]�y����>�6�hF���ф�(��  ��� �}�hEA�� ��z�{[�˰�6��D]�m���/�/����M�����x���K��i�������ʈI8^t9��%�upmcS�k�ĻW<»�����ߟ�!����O�!P>Ȯ�(v�G��{sG����G��U������'T8o�>�W"�z-X�A^�!�Gڃx�hN���ة��o����г݀0ͼ��r��T�q:3��e.�e�J_��*�7�NN��U��5��/D�qx�-m�����.�w��@��C�{��ۜ��ѧ�/I�s�c���K`� s���N��*���K��U����k���E��
|�$��������y���1���Ƭ����VG��F)L������/+��
nї٪�dq˘�9sd5�+�՛�䔍z%b���0폄�7�=w�)����G�pH��Re@�*��V�Z��͑����[���g�4:,�,��K�7���-��Ѧo`�o��	b��KM��f�X�
?���QPm�9a`F>#4{;���9x��bA�C��S��o\J��zs,|���=���7�5��7N�
�̈́�I�w��f���]پ>��Qzr�<��霌Sȉ��ect�"�X��Ɨ �qy�?�d�M���D�І�
ޜ���l���W+4Ӳ�j�����ng�O�i�v=`�W�����{�垼�����0�����g�@��-]��Y�On�T�P׏�X��WWb��F�u2��7nK{��+j��e����z�\V�
F�Msk��d8�h�S��Q�f��?,B��<
8���n� p��ǥ�G ��i��"�G����/So��z|!4as��0>�9���Lc�������
�QP[�7��:M��^�,)rG��������<ܳ�I�FH�,�]��ח�lm�E#W�Ƽ	0W��n"Q�{6YE4�Z�/|&��u4z����<����>B�a���u�T���+�]P?d[�>|*�n��V%^D�(VM`-eB��mC�0�;;޽�NC+�u��P�`h�-�{zEQs�k�^D�O,`a��u�/����g��0� D#��Ƿ˦�����d����<��:�kky4�1v������~����{*��U--}
nⴅ�U�-�w��r�Y�Ié��Ėe��h��\젎'm���g�q�u��]?���9�g�ݶ��t݀�g8ռ3��Y��;t
��]p# P`+I[������\n�0���l����!Ԭ��O�`"��D�g ���צXu��ܑ>��??^xo��UӮ�oP��lE,3FMA����d�FUt�ɇw�Y���*��^��`��ㄌ�;S�K��_-zۼ���Y<e���t�9��)B��)�m�TD r_���aŎ2Zs ����*
LvPМ@]��c��b5#܍����@��X;�����ҳ�;׉~��9�Z�1�T�u�g(`����:�Tv��9?�[�ޮ���.f-�	է(��z����<�=�T!�=ҖB���N3�+eo�$���[x����mnxr8ٺ���N�tڸ���%d��w�hp"K�W>;�D0�:��p'y!ŗi��nsKh�����9�R8C?���C�.N�yh����H��Wf��(��S�#�l\��EF`��Ue+t��pu�ѕ�0��~�:��������m��6�P���=���`]��z� vn��k�9?�0}�����k	��d�W��n�ͫe&Ĕ{��ᑟ�֚|CK���$���%9�P�h��,���oo�HEAo����L_ܟ���8I�dt�fGB3onK�Y'y�N��t7Q���gE�o�hR�R��8C|���0�=����C˾q	A���1s<1�U�I����2����7�(=s����'��6.��D��(�62��|v5�v��h��އ�X���Z�/�B��5��; ��v_E�U2��{J(6b A� �	)OO.����|5BL��)�#el�*�J���/vJU-X�aڗ�3�W��ي��T��mT�?P��̞+�:�"�"I-F��1N��&8z��5ʈ����$����m�Q5Bۅ�􍥸s���ㄱ.�CG��B:2���Ǌ]痜Ⅻp�nH��@����\MG-����I?�_��B2��6(%�Ē��a?Sm���h��H�xV��@�۳SL��ŏ�ң}]6�e�0���Ⱥ:���je��U<���������#� �����~bt-�<���(vd�V4����g� 3j6"Â�`3����/�2�t�41��.s!k��jI Em�~�ͧ�b�6�
ߕ���� �>p������Wջw���~�V�%���U�C�\!�a�E���UFy�Yc�|���K>Ջ�)�{i��u� =/�T;�[��}D�lt��X̀�A�Oe���))�ug��/��V� ��	��ƕ>Y���x�Q&�3q�>$��g��
z^�9$[ybA�P��k�m�SY��l�"�'�	�Ffj����^;��d�G���)�����X��+�>rnD�3�`#Ւ�@CAj�D�kNw[ş�6�~��}VG��i�}��x�\���V�g����:k��ĺzVE���׈��J�͹���}~�Z �E��3vg�u�r��.�k�v_�-��)���܍�ư��2��p�s�n:A��z�� C��ı�Y�[��:r$=������?ԋL�U��oG_;�X�'҇���2�@�t���^���p���`Uu�Ќk���y�[���E,�\G���z�}A��FT�YC�٣Q�Ja�[~.�z�3<�m�	rL(Z?I�&r�L�S���+�EGQ�ߌ�/乥�]���7�Vӄq���v��.i�f!+�%��E�}�?��Aa�&n9<3Y|�{9�"��Y�q'�Է� %�S���	�K~��0������.=b�G�o���P�$Ӥ9V�`�ፂ2Č�:�(�">Fv0T������N[D�^� _iv�,SK��L��cz�ӊ���a/����p�e����3,\<���?bQ��b}�j�$�����gM����3�����3�"�Z��~�@:k���z���8fC����Y5T)���cE{zRphi�I�	1�������+��E�=ʵ�Q+��8z��ן��c<� ]�{��+w��c�0�H-�>9HR�2�U�F���z{dA��.1tu
��¬]�.7d����F�!\"I�qF9�)^�<�hÚ�+�gb\`N�X� <�vex��73�q����Q�w,�EL�V��rWk�#!�4�
�܊���Ҿ6�/f��aJ�ځX��?S�H����f0��
�%�v����1<w���	*��
o�]��R[������[��c���"N%^� ���ҟ�|�;��S����9����9ϱ7$a݄v���z3�{�"�2Et'���*l��TP����q��,�F�uc�PE�j7��6IC@�N�G�5uI����y�gUJ���pn�$XY��:�.�Y��L��/~��DYק�D�Rrz;�i��+�����em�{ō��2����	�w��ӏƲv�a=������_��` `��.!�I�1�!_�	�ؕ]�P)�	�Yu���$�k��!\�ޑ!Z��Ъ/C�5˂�ж4ܭ����Q�T�36.���=��X7Ȼ��"ޫځ;c�b����K=�f���c�O��	���<w ƽT�puA߿փV�:��=AІ�f��T�56p�$���*��%���|!ج? ӆ��T�ļ�O0��D�����h��<�3�����2"��s�U[.d+�s�-(S\4��p]+4����D���
h>c���@5d�_D�.j�vN�Vd�������
g�=�J�����u*s���	3�;V�|:�F��3��){����6aϝ��E��	L�2%�{<��B��Pm�s��a^o5�\����#�M�C�j��k��\���QC��Z���{N�3�{�N]�5��^���rZ�(����[1���ޓ@MB�7-I@�k�
'�����Y�*9E���]X�����q'��L�6*����\�A'`��3C��hT�i��r�30x�W�_Tx�N7�N�3���&C<�Zд������CY2[�K�:93iuGEGa}����h�k��Z�W�'���Ě��� ��L���k�0�G�m.���;��Wl�,�w��O+��~ö:cJy@���dX]f������ (�}B�r!lU!x��l?�s\��t|�_����ȩY���o�գ��j�b
� �}Sz����k����e�����q2T֚2	 �l�̶�>!�]$������jR�4Tu�7��\D���MF�9���r^��=�z��S\c�>�,��X��(VP�(�;�E���M����<@ķ��8�7��pb��lil(��0����m��:��U�G{r�ŝ(�����`�-<��D�E���߳�����h�d�g1������$�d|璬�LJ�KbڗD@���!�^

���|c�OhM�#�[��|������*�Z���Al�B���$&��h�B����:G+&����Eİ�@Q�ꏢ�`�J�2�e�	FrS�1Q�p�R���;2p�傽ۖi8D+�=F�]y�?�:I�PUK"�W�B���"�_pN�G��*b�!�:i�:`7��]�`�[�3G��=K��y�P%uO��8����F˕i )%}�8��!?��䭡.LX�]�e�}LyА�������p�)��7T0L-r�K2p�y�oݍ�$��{�C��6:�-�zȾ:������߈3�1���Tf}�����\pF��Ä��j�.ex h	�W��U1[�r�h���'�!}d7�4��iM���/���A�	�y�d�n2�#|ӗYC��hђ�N+�f��� �P����r���掠�
Sd'�Y��5���+2{A��o���s5�CA�m��M�u�`��He��z�r�R_�=ϥ,�׉�T]k�+ĵ����:;Yt�%5����FV���ZG�pôV?[.�!��
�2����Y���s���j�y�`�C�%������Y_�Ό�􋔋G{��%̘41Z|Knp�P	DO*d&u�#r)��'�C�S�u���s?���&X4����thM��]qZs�-AP�]������j�Ƹ���La'�*��a��k@��6Z�vQ�u���&�'��UGe�=��N��F�j�e�B�R�^�G��ũ��;#�ï}�Dv`:�{P ���Q�2��ȥY�+�PiQT��qA�g}!N~1���:%W�[�����g9�Y�9^{����"�F]3���-�vW��(������g�,�I{���z\ B�I)_x��h[����-6	��i�d�,�bjt�������1g�SH�L�d\F�d W��$�ka^@��c_U���I�������a���ߪ�J����L 1���e�y�0��%8�������Ғ{1��!�X>��j�5%�ۀ�|5�
��^��?�s��w��|�y����hY�w?¤e.�(B�(5�G���Ĩ���>g���ox��(۾7��фF��$D����Rf\i�lM�7x��!ݳ$���2����+�Ȉ\��B�?��r��<��Dx��-��D��m��[*���ޟ4p�M�F�O�78�Xۊvg�J�UĬ1�F�F�iv;��+�@(�b����B&+%�W [ѾW���>��T�M�i�^!-z�c
x�ұI��+&^�+IEg���Q]x��rzlO��xhq�!�9W68yB[�	���}p��qb�'"�[a��~`�s랔|�c����,"�2}q��9�9� ��R6�����$
��z~{��t�*�O��L�2ìD�k.<@�[J'�#'/�](W:���ts����M�e�i�E@�|��?yiGc�h;a2�E�oQ��!`T����Žy�ܹ���"c��7[��H��>���u�"l�r���Îa,A�)�H�G��3?:6��Z����L;���Q�G0W���:L��E�A~��_	�$�g��V8��gq��u��XI�K�����e�	>[�o�N�j�d�T�t�D"�9T$�jP0��k��z[�<sW�ءG�ǋ���x,�N�%P�B�U,�	��4�ӧ���
��s~P����[$a�\���>vc@M6���%���y�*�1�`�3J����\���jX��Si]zu 3�Fj�d]�U�~���wj������2����1�Nfm�z���h�=�W%s��ӺG�:��a2lEo���H� ����_ؐ��Vh�%��w���L�g�R�V(o�4^�+��	� �����	`���c�q��i��������}���7�p��m��y�Bd�0�Н3�:�*��a͏�E韮��.�wY�S��.������Cݕ�G!�`� ���+FYԮ�}�P�x�s�a�1�]ߜ�(��g��[�"�FSGQԀ4��i����	V[x��x5?Zy\��@R��Gq�}���(#!!x0.��'F���'8�$;�M������i�$�'�,���A�z	nVѳ�F2}V����'mM>[��jĭ�_[Y)��|�a���!���9=p����G����@�	�.�N�������Z1l����k�)ɟ��N	~��u�O��@�	�� N�������0����TO�9�<�H(��":�Ip�0Ѝȅ6 ���z��S!i# ����-ТZ2p�T��\&�H5��%����*��h��1��x��R���N���53������18�o�	�Ď�vo�+ͼ@m��b�7v'����cw���#h�i%#|�����R�\�݆00�W%x���`�2m
:�
Di(5�9�v��ܡ���Fsm�0)u�S�����T_����~~���td�[sn�E-��ݡ���I��^7���Ka#�)�*3F-,�b�ǻ�|�0�H��ұ��R��"V��ob��?��LMm�9j��,��"Y-a��qYI��K���|�����N�r0��CFzQ�l���|$=�>qI�aP5	����z�/C�>\V�1�G�q���);[yHTe�Y��O����r��0���MF;<�į�Bغ�:tθal;G*��yX���s:Nq!N,�N�k��v�6�T��E8
?8%pyߺ��>fs�RI#2aߦW.���V����ۤ}>�9%	��� Xz�)��������U�L9�[���b-�E�l�bd��9��T�B��P�����`�=�-bX����Y�ѧ�Ez�l� �;R�XU_H��y�����w�<]�`	l���?Z�W�9�{�z�j_�"]�������{�q�R�%V*73^	���dܷ�>��=n��+�.X�vf�e 7{�-0L����r�f["Z,�$|��P�0En�� ����ΙU�Oտ)H6������K~庡���=r*�z`%�����Npu=ƕ&������Fx~��]l��.4$u����F�W�p���Bm�87�[%�e���!���^�����4���_��mTix�R����C�\