��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,G�ss>ʂ�C��S��D/��mD��J���Y(�H���U��B��Z���qw0�Kǿ�(�yvE�e���e"k�^C	��?��*�#tZ�����][�5�zA�o����	�����^L�F��A�g=��М��<_C[/�
�̉2^�����|��ȿ�i�}��=,z�%\�HA&����>=��O�t�>�b�IN#2����x9�̾����H,J:4�ld5�'�	�9#�$�喠�P�I�%}�S`);r䗞x��Ԩ��^S�_cw ��?(	H
�Q8P@Ϻ����I%���5U3Y�o_�';K��8f���Gyw���;ЦQ��-#)����E_9�C���z;�v�.�q�]����Z��	����GF���?�Ȁ�MG��^]�j�k���8?.�M��?�[W���j�k��Qa���5�#�[�.��SH%��l�,̚`ſd���?ψ�b��r^����R�Ϥ���[���gW���ǰ��uNv};ǳ9ཀȃ��T�C3�$8���ǡ6e��m�<YT�X3o8�WyQ��r����"���t���<v�]�q�)=�ʳ���،����u�/Q��r{��~4�����%�Fh��7���"�-��_o2�,M�� O&|O
9�g����mj�{�
�y"�w�2n��vJc�ȥ�x��I6uZ��L���za�$�[n8�vgRˮ����G�#���?3��y��}s�	n�i��_5'^�b����]&�k�j��*{<��)�Y�����1��מ�۟5ݼ�˖J�e�dJ�}X10DQ�B�n��>((-��st�8qDH�v	�IcBXiq8�>�b��
MG��=L�W@
�$��r�p��t�d|9��5fj�Ϣ�E����z�΍�"ͯl�=���]TV'�CF�����X�8T2tO]=fN���3�)D�X%�	�9Pck��X�Xa7 2�?�k*=�UcP�9Fe՜U{���*w�BdĊM�D$�K�l�i�_"���� ���z��=�uHg�IT]�Gdolʵxю�np�d�U�f�gv���������}S�����I�:������!;��8�r��j�"t�+U�^϶.'���D`�B`Sx������J����s�����ԣfǧ,�������t���N��qm[�gK[�S\����3�x���-�w���~ձ�vi.�d,�����/��j���J��0�G[�w6��,J��6��ь�)�k7��C4�a j
����_�RN�U��ڛ�b:;֠�?e���x܄N���(�q�T����4g�:���<%4�B����Iz�׍���@���'7�A|�&���Ζi��c�V�{s��x~}�L2�@츣%�	��ֵ��Z�����������~�3Y-C���5�z(K��r`��Wb*Z&��5�g=��v�$�?0�^SE�']�d'��-#������+L���'���D39��^Y�}P�2x���9���*��wLΣ�YV��~�<��}5�Rǫ�c�d������s[V�22Ffτ��Qs΍�!�������B�X����� x-m�u�V_�m��6�%,��݂�-�-�nF-��H¡�x����,'@yHĒ����2�A|�
��'Ek_�5�:Gxӊ���Vp�#?J�(-�FF�� ��l�]���é�k� i��j��4����-��P=�����DmU�)����F@��wYg	i8��_Q:�_ީ���5օ�NMO"��**��(8�T�duA ��f��$tgA��?N^��B���UUZ�)�8��n�3������B����`����l���R[ߠ{�D׷^YhܘX���zP)�d6y�����x+�,���bjk��e���E;���Q2
�TM�_2�j{�,T��OQ:N�6�3lh�C��ǚrT�]��/���B�tu`�t,�����dh�ļ�����~�r��\xI�'������_����b>wv�q\��t#�4�+�xN��d|���4Aɔ��NEy��٩r���H�Ch	3���	>͒�* ���#�˗�k�ZM= �Qp�/����G@So�)"!:��?�L�]���-��"ؖ�K�ȼ�c�x{3+��Mδ�似N��*a��(��m���/=c�%B��)��o�c����}Zz�-6j|DWT�u��?��O�\b�j ��M�h���۬�j�U�� ���[g.���r~q�����T���'�[���i�ڗ���fM���P�J5��H�g8x�'���!Ҧdd|�ϔ������}B�;��AR�N�0F���t&>�1n��͔1�nI�pj@d���s� UpH�aףx�8�?��9\'dsI ;8SpVGu�s*�/^��aq}]����
�މ��l�8��v����m��=X�<��u���	U��[&.Pxo��*��݆�.��44c�l�ܐ�$ff��)ν���o�u�K�ȷ�� l�g��y����i���E�]~ş�r��ϱ�I�o����Ũ���|�����ǫ�/�� !J���I����4-e��,�d�#>v~��/Kj&�����ya�<��$��I`���4g�{as��n�Q꓉���^c��eFY��rȤ����#�����p�w3^�s�
T�,;���N�%m�[��&mv�;v���]�s�\.;�*}���L�ڂ��}�&��.��%��c�MT��c�_\��W;��(Vn��pI�q��$
gʨ�\���)d��� �{�:���!;������:$Kͦvfs43�#���=�h4��L`�I6��h�>���L�G��Nx�N��wǫ�GQ,�U���c�Ѿ���s.f�ڤR�t�����Ӿ�����CN����.�U�8��hOt��S@?�%,9!f�)��7�~a��^�����9��/��-?yY[�ӝ|����+ �!����W��H	}�q�W�_��M�{H���u�k�	r���*>vI�8�$$c�t�jIN�q[�."�(!����d%�0lBӪ<����Iff_HH��;l�s�G{���{�������$X�2$l��H��!�������(�Ԅ�駇b������9��g�_F�ށ��470v$3����L��?i�(��UB��(��|�ީ��%m���x ��Lu�����D1C��&����OA;�7S<��]Y�@Z�C�����(hW�P�$�7���+�4�!�'�-N5�[�=�%]���Zr�Z���ƻI<I�s�4�-�� �)	��[��$�Y�kй5�ӘY������K����M(Ze�۬���PbΛR��FB9�
����ˇ����l��'��-��^�8y���T"���Q�1!7O�Q� �Re��]rD���T���H�h�Z�4Y�i���bs�ȏҾ��Z)	�9���)w+��vR���E��J��8�t���=���D��Q���eh������C�>��a�VR����x�������m���٣Ծ�\�o	��-A���\��A~Llŋ�b��Ϭ�3���(­eH���t�+�gl�u_.�E�B�ά�Gh&U�_���Vt�2AJ�w���>. ;]2v��z�W���[	1���.���j�6D1�H��v�z�B�vu� nk,�k�bY�)����C$N;�d_c��3o�#,I�ZC�{�=l2���\�q8��K\k��y����2�!إ&�L2�}�P7���|T�K����)'�X�^�J�tJ�ޣObFRh��bd�Nq���f�uy�G���b��������X�y��>4Є�����M�n�I�2F�d@��sYX���Z�Q�H�@�@��)�CQ�k������D ���vb=:	�%��l!ʕ@-��l�f-��WҜ��^r��*�F�c��d�ªX�ɒv����mĘ�)κ�0x3��Z�+���j/�L.����I��I3�{�_o�"az@۸�t�ɟ���ORJ��n�5��M� �O��*QX�I��s&s� �O`��)�&��:܀9�_�rb�d�:c��u[���R�2_M�FW�"p�^�w3b���l���b"櫯Ĭ6H3�|� �Q�v�	�k%z���6�Ø��_xzb��j&���D����L�EІ �U�����$�|��)%�K�i���v�J������e��j蕳��i���@#>]#1����u��4���>�&OPO�g؍�G{�q�N�GVFC�<��:�m��q��vVs �2d���������ַ��0��*��3Ky>P-f��G{���مS:Z��j�M^�&��o��x�6�n���>w����H�n%x�|�S� ��s'���iFL�bN�Zu����RZ�>������]b�(��:ح	�����Mե�@�D�,�N\�s�ɧ� Ck\]Gp�V{���㳤&�=SmQ��	�(tQu����Q�6.m�#�]������M���P�X��#~�vײr6���.@��D�-cK���ǑMǸ4�^;��<%'�薎���l�����!�.��-a�s�u}d�Qh�bKM�ۏ �Az ؓ�(�u��%������m!��g�� � H�H$�ŋ�6<m�2����Qh�YײN�%��vY[��k��b/��*.�h��Ҷ�KX�H�5���!V�5���1�%R�]oCg����k��T�6/ӹB�Q7T��7}����as�>Ep1q���j��ŁdL|�M�H�S�G��y��%E�a�'�y��黈~j/ӽn��Q�Đ01wwي{�tp�^�m,�µ&�����.�+��D��'��7-ǧ9s��1N����Z���d�C��3p:/Z��n������*�P�XL4*���n+]��րP'K`\�|>x�j��>�\}MRwˇ�G�"t��d竳|�7�݅yJ�;c6�:Z�3��'�5&u�ǧ�ҍ)���=�~A���Q���}FҤ�X:dۣ.��[�I���x��J@h5����(���Վ����&Ɓ�]2{	e�r���@��(V��V�:�4D�\vw�W\����Z�q�D��/}D���9���o�tǬ\��Bk(�b��%OGk�D���VbA�Z�@j
�8������	���q]l/HCy*�n����ٖɻѠ%Z� �j6�	�*�O/`Ѻ�P�I��2���[�&�|�=�e�N����$r?�S#������diޛv`	�3�HI�K��M�E��"�Ő����]�o� ̴B��^ �c����.�w��K�œH^����;*s�Uhκ` E���Jr��I�g5�e�B�a���e5d�M��>jS�vJ�+1�ڗ��y܍�-��qf~tuª�#�����s�0]f��N�Ci�tw�<�VV,��O��Z�*Yy��*[�I�����%{�n^��T-#���)�lܷ�,��,��k��Y�)L��u�;}��9��PkL&7hQ<-��m=�*A�yc��tu����B>dk��9gZ��w�+�p � �3�jN�6?�e���� t�=����6iA�6w�}y���މ,00�j(����}�2H���XA��7�栴ݬo+=�p�Q�z�Dt(�{ ��YJF��������6�P��^�!�r.6�@C����OGU�&���.?�Wれ�?�٥����e���V������)j��J���QOe�8I�����.���{[vY��#�'���%K�Q�?��]D����=�__�
`������͢�e^N4YI���*�l&1L 8M"F>����8>�%nJU�B_�Y;�4����L�Y�J��N�՞�y{�����8��e@m%s� +y��C�4_��V�7�i�7����̯t1i���_��IW�P�Y���r�L�np �!P�g�A�S�'�aU��K�=���Ĺ����_���2�`o�GKF��I�sOdKL��[�H���8�$|)�RKh!��!�kc��B�٠�cb�����_V �/��<�Xz��D�<�#��"�A
pn���y��'��	��|m3�Q1��D��n_�Nj�!��y�S[[���.��#�\%�H����z�ٚ&�@Kz��fNR`���L�jV,�oI}��-�7X<fZE]kl��)������F���sw�ZݗK�ٍ)��X����Q��#����F�d`�e\�) 3��
�߈]tpcz��Źr����=UD�[�!��EH�=���ZҚ#��^�b�$*���Z�b^ȭyn�����\ �ts�߳ĸ��ZU�P麇7[}�c7����LԢ��G��ߋ��Yv���$�+����d�/�I�7|G^g+�,�	XeΆDg�K=��~N#��	��8��Ӭ#��˶�:��,b ^0r�Y��k�N�;+�(��&[@�.��E	T�f��4i�D���,�M��͸�^�FTf��K�"���)��ń�
�0��Ĝy��q�r�S��Eo�D�HM�x��)56:�%X�}hMSڭ���'<HlB��<���l{����uN	���:#����jg9>|6r�S�>�؋o�O;�7?�ήn�AX��{i&M�$H���b���a���7A��IAT�P�k|�Pv��0s����6j�