-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
v7dFfoTrOVYpsuW34fdnyJGgNtxF2Hu9SpzgQBVeEs8u0ptEvmUDNyyHlcghLTar+tx0XOana/sF
gfIhw1ZSvPHk9Pm4UQcLV28i/6EQxLraK12uClgiOLRP0gxC3+eiu3key3+25dPVmcaAtPSZR/O3
/RdIC3VtpXgwbhivLBICNv2PUAWrs/vYwqKdtDa2VTe/YptKXRMJ0nLAqhXTYoM7TWGeDS31F1PC
dWj6Pz0+udZBSouNMpY3cCu3LtYucei2y7F0FBIueQfgcVI1su/NP6UqVvWXNlHYP5oUyAGa1UzF
EPfIJvEVu5QWqPyig1C08E4oY0wdhKo8874nYQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 23808)
`protect data_block
9wgVkyNfNmNxmyyt4XqdHZIkxsmokN/HI3gMuBzAFAXiYXDOZ8QlouqQRaFG769uHpRnz/sxEn/o
y0IBi1QRx7FvAwHQA4S6qeYFzo0D7xNCz3OpQhWbKwcZugadfnFMrpiu0yiPXG9F2totHXe8/aqF
iSKvu0+W7cNuwmqKC2uJcbb9kDfdusIWOT7t4LuOAOLJaWXEZBzBlMbe8sE9/BFWFmPtcvq7ql+Y
AWxYoWhtKX9tpARIhwN/pJKUD/nWgCSIAOPQuAF3D9Din3uPfm2Bp7N1zexoPqz3bSO1ft1MNJal
0ODJVK9cGn8W62PM9Cw1hSuAFfwPkZre5AsYsNSTVOF282oV7bACR/1/oHoiOF3kv3Vjrh1qksji
g8HO9fXxfvVOMaWhFXGOEjKOby+U6JN3OGBEbF6Hti44JIC7jl5Z3EVBYhODQMU9GM5Omx52eodM
wHK3s0IBGL+HBbCAE8T7fdhexH/H91ZYL889vfZe2HvepbL55vKUOMPfzhM0Mwc1q/Whkee3+x2W
0WQxnZSg7mTZWUN0delJS6XZAqRV7PARC0PRc6CL9yupC8Q7RHFfotor3hHkkpSTG4l/m4WnNHn3
Tuu6Gr2pW/rIwEFA2e3ZvDHmTFcvyQgTbhMp7W9Gluc32mC7kK6MQPYaTBfjsWcgyBT2O9ueNUMz
FyTKN7cvmZlRZVuEQ4MKvbNC7eLeZr1kbwz4MJhm1Wx3afFnNuoSz6g7E57icoynDFc6/9Btb22o
r/ghLHdI0mhawSxLmZeJvNhz6fIhoFIfexMC4cMh//oLhSBGk3ttqaAteKelq6EUt9wPDCUKPfkw
/5fr2YbGG+IVO5X0iYgyz+GRGdV/eCmFGU+hhhoIeWoHx7WHgeL6efhN93tuVMGTmXGzfe8agcNW
sybAlXbXIB9nEfrspf8qXVR3Ck5AsZK0zDASuI5oi/S0iEPa//Dn74FkaSFBe+cDpSTNtDevBVWp
n2XaYhYFssIc2T3pgVg0yPsIHBf14ii6fPrWQT3OA/27L7nC4d4YWVO1MbpsQTFcUPAzcIgwEAFL
nkXyck0+Q/q0GjMmSwWGZndOcARwqKD4/dV/07hHhALdySsq1y7iK6x1NkQDEhaSInrrEQg7bdw1
j6rAK0v86ez6zhyPQrLjQny/cEXU0uOxvn+HAAQ9xeBozN3HzmDSWaxk/DAlgDrouQDThbkBPZNt
BXFIlYhU4E5C8Qb4My8pXmErRzHwVJBUfpvwfZHXi6BjB3tRfBGyMTnqelU1G133eE5HgWYznUKy
WLawZJG3zW1zKrJmwvJSsuLo8T7IjAYDCKYLb+w4lQMDzTGJs0gjV5sUT4XGqvJDMoNUD9EgWONv
EopehrPt2YBwX4Ynzm7CQWI1JhpUr7q/vhAbxkd7jEyMIZqNMJBQTzeKtpk15J7nPKvqVC/GfJiD
AU/eLdb29Y6XEMwczPyzpr58IaPr9lpvWIFej22gmdkCD18dKvstpkjnuY9mXoW4G6F1KDyC4my8
fojH2m/ljA2+m9IjC5gVI3K4HUfzcPzSiyw79GN3AO2mcnu1nYAvEjHIe6YwjF1OEEei+dwiDV+k
SCYM80JpIUNTHiyw/iB8SYdnAR8wMjKXgafMS8I7pD9GyjEWgm5Jdm7QV6EBUMa5deyfvQ4oySsS
+IMZWYRLWw+P0EzbjFcmthJU86zu4No8kU8PRIiWWwg7C6HGzO5O5r6MowKdB/H4NcNH28JnTCmX
k5auWSi+ftZM1tA3Bh+lzqHnYuTyofY+irdaQLTaoU/5jSXX1VLrgDRuKBJ2w4mchhwee9wOIqDt
pOv89hDKy6CMOL8nNiPR6NZ4jtsWtVZOsc0xDKeIsZB6r1bUoih3kjRtRXPDlWy6SRYpRo8glrLp
wJDqhr3rhHy8haQFhuPeU1paAPAV5Mrxl00ITPx108pqWhM+1IHNIWgC2bLk3SEB7SD4LjOj+TMA
hIS53ixX198u8zQhNdLjHrYBkXg3ZF2e6qCVnA82M8BPtvfqK+E077rycIIfc+ncu/OwrSRoYywv
5DcxWN2vtpvQYmlc53K2ikCK2J2dSu9LWTl3zHaVZzuKJq3DdpmJHjiS49mj4RR+S3I4RvXfxkDP
YIz5kl9cBXEQRy42J3Q4NsHt5CaAWQrDJE7o+OoDZLJf/5PSuQWm6jhS3qLPLMxSsjvidxNzY8r8
9mEuluHGKdbuaK0Jz3xifpmIj36dSYOzCMUlmn0wJ9RpZFpbOzPrctJHKMzr0xMquTfZlVAvaQh8
vU/F1bwnhcvLFEV2hOnz4T48XiqhzyHby7voKm73AV5OpKDiB6s8YOIiZcGMz74bWhS6l/T3tMb4
q6bbkEBIuAjWB+G6wx77f9MupDbBQZ7IZ4HmhB1uuzRmFAnwdXQxflpxUdNdPboczifa7BrthC0f
m/W+BIKSkBFiJJMPs8mc0gq81RqVa8QteATShWS6JOzKgX2yDIPyRAtNKA7799nii1i5b6//YPuC
NmEMgUvP247oVhToUzrJzgqqGv97vNkca1t7vlOTX6Jb2zgcLRb1BIylScquuqmyg7mMxA/0J6u6
714uUI8clV10red4EcOy0qxf4SW8ro7RiowF8Ib67joPYEZtkOy2HKEVxHy+9PXfsFCSy5lwpWwE
fej7eSqVnW02qIHGYu1NBYfg2UtA6V/i9olH5gvH9s/t/QYtd7E8u8nsu+DtFCB7NhpCh4DYcTt5
r0cPJxXxkatyx86JWn4XGuHWQObjF2AGlGQzFRlpraRQKyiJ85AZ1DJC2+nbtO1t/hXND69Kru6L
QnvxrIoCYPDX+iC/6WZ0oBxtwu9Te5iqGNS+JSTse+chHJFVQ2MO15I7SxbooJqO7FMnEPycklFK
Gpe+9ZPopRzYCqsda3l325DNLZNmN1yEaQsQR4edE5punU1LXEVQF2h3TpyFCDWvC/3wCeSOTzKS
eGX1RH4QzWNHh/Q0U97Ujt8q65cDS7AzkYcefWqMQEt9T/iN9bbBqYBAviNiTiNaJtdJfDhsAL2B
VTS5a31HbsviVfg0laa6Hu/3PFKk+j7PS3CSVq2c9FTn8o5AWJmA6V9ged3cl39X/voNwwy+e52O
2755axM1Bq8ssEzFpjWYQOZ6n2Gufvwess1GrmLFh1Y3pGdrmecTMiumfqcb0eeshTEO9rEn3GRr
3bIj/cQWnfbTzaMYGY5+p+wOvBX1PKCY3/H9iVIzTWvQa8O+twzpwdWlMlryJNVqs1vKpEIAk0Jd
TNe7AAd0Sdq+mYZc6kJhngUPrWXaBxKV+7Qvn71Ci3YZbArdDZ0CO9s6tHdCSu0VMyVze1IoLIpl
KSJ358DgB9LiLuZ9JT8LHmQdKL+QLgVuwxUBCRlrkNGU5cgrllFL8uOx/c9S30rjMW64AjT46DWv
z+xIoXo/+F0apL/8F00PKzfC41sIV2iaY062VTAzM1eh7HfJDk9Ql9m8oX7YfnWYVQ9g3NMWvwh5
s5yRtVovgxYbuMYvTcSSGbBJoCNMS/EonSt9MwMmbNkeOcfH5we9zC9qRMOUrHMiwxh6Iz4GNgQI
ry+y07Dt/vhozzVL0hY1hwBy/2cnWRhNzQQcwLlwwlClpyKR2WYBd21FcbXS9Egtv0YUkTAafqpw
cEaJm5LKKjrsF7YjGSSi8HtND1XzELb8EE/n/nujQWSjM2qXcf/7E8aF1JRZCOWWTm6Y0+YORTiv
1oSocbUhokt22ddY0c67Cl1cPLjTJYWrEnN9leWRK6H22rx/0voPHOrJglQpO/4HqClIOqp7etBN
zTzvZXJeGLNLNiXhp4wv/uxvk9oPeWTrMfrY0ZEDpAo9PWKXBPwmo9252Vk8lsy6eDGgzwVZjgU9
VFbp4R8Iq2zO/1i77F1CL70Q++7xE69U4TysgsHcbHmBjrQy2GI75jTthVsJYg+dR7OdNGZzJIzz
DzWcTCXeLrilqflf2eU3XIrgftJZcKP83z5W6YzmtK6zoAsvv+2MKFEG2IorKKI1wGn9Bmf7qStq
rWNasAJQOrYB9smP3/QkKeJDmY8rq+sVaVwv2B8CAgKJjZK8KlbMH4VuAtWS3OKk9gS2MnBcRbkY
okei34Txdh+sKO6W1PK5NqiCUbsAwWdX1dE7fa6fxjHadS4J0TQcCwjR8sagGjLG2UbTl3V4+UjU
NUl2KGrVLIXgGeBtlzBQiSxW8qxtXNIXcMRCOzQUTRMzznHwA2T0FC+32l2y2SvMh3ZxkykyWZIw
Nig7nt+2blibwUkDUMdUjfH9MxtQQ4GX1mE7RfhVvD4iLMOsDyXlg6vf730Fq8QTcZD1Aq/dXmpx
OfD+fUu0TBQN3zO1sTQyM00gXeANkA8avtfAkeSZ6/w5nX22q+q+nIL2aSQoo2SJknyx2KyKpbRT
6dPaO3nN/NLB7kcPvvaMrH6DY9WeZjqUp7rijJ8Nro0d8jQkzHHUpGHn41kdggYvdVs46kK0s6cV
BokHKoONE7OT54IxgfYw8taUlVtqyDXW3RqWExGSPVsDTix5MBmbQ5qNQxpmr7MaJ95H6aUZk0Lk
tbmcpsno+FT0Q5ntyV1zhXFrmCzDvRa1bdmR1RtDUfC9AlVO4cXpFcjzQTbHirgc+VdEUwO2FPki
ImGNU0Dy9g/BKLDVaNm3du0x/kaU6GiB1iJDoFyfRJruZvPFtlqboCk4y903PuC0VqH8i/69NYYa
AjeQglowkoNzvZeSlgrlvdbLPCorctqurnVghTb0Bxb3axWyOiI5ogsuqYwVAf1FLePsQpitYTZx
VekkanQWBl4297aJHMPabicZccqpWJagJKmojUg5PNtDDoMpRxWtbdu+cKBHiopoFwsQNnhFXocd
wXYw1BEWIHLsOnCxuFPz5VEIyd+2robr2KpyFNuqEut8J0BqzaXB6m0drgOtfSViP50ETPYY19pI
4RObkaSmhlbp3/yvSt/8KWI2Uxoshe1UoIM4iEAejVUF7wzbsdaogjiiupqHb6/6XM0UnfLFrZPd
kfwbUs3+fuOFAYPE6/EvrhHRvqIKhWt3l1Ac+JfFGCetRyuS/82Cjh7/qStix4OVNWl6pLU1Le3x
9X9glIK5dWwNgF8s+r0o5XYPgOVeVKzQpBR3PjBOZeENx8ZXFfBjMzBuHu1i36UP8pG4BfKXNe8D
FpgHPNYBR7dWsVVBrqsEEMxgbpItU7Qvfb84xUQsNrD9d5QzgG7JVhMA93YXhCjooqVhqIygZAmb
cfFqH7RIUL4gvE0aNggodW/u5BnhUzf0YoMDdnr1GJUcSXy1zAWlYF5ETmhRhj/ZxmvZhSLlmr6l
+WWN9fc8YExmeVTCphZcOz4DOMkPltmnMzkNqQn7x2yscmliC+PvDyxfAl57HG4oYJEBM7MIYUzj
LtlaIoFjFbfz/ov7XGXZ5/+j1HFbQMelsZaJAhGSRh/EqvHHaHGKFoJ+pLzwr3ZxxGZMbCm8jsBD
pLU/nfkPoEnWfV3a0eWkH/6R6oeKStjb4R98gfWgZlAsley8EE5W1Z+82HkTQGjIBsd6HaETXD+e
gYlPk4ApZgi/Agx322JE/iGjyO7iPkoqTnnOtTzSkMgTynzuKC1vxhPDRe15EbqYWd53pdqgOs2I
vaNNYikHXz7ou3jS2lHxGbcSYMcj2cmZOOPkNFU7IjRexH7imR5YxUfvCMvPk/pJU4vyqqiKvg0Y
xlkkwjCziH5203OqzRmlBqGhTuiIqR2bw5yTSm/vXbbCGAUMf3rrGy6+UUQuEnKbBDYRlF3JR48I
8unL9MNnfrxzoxKlHipu+9ktl9SN7cekcDuJMD0ifmjIykLMUCy1CPXtZrwWrXtbo3qm8OtPBqrT
DQ82vgOsk6ecS49rl5ykAIhNmqiXlpiQJi0sWqyvwWkByqNMjDwOJh7L6ohEy/PQU9L9SVS+vx4E
L+DIQEunGMVpk0d/roUJM0aUXhk1BECdJK78NsExPww7wPy/tOEj6FxEHxkGTLdQ26iC+ACNYdYR
Mv0CQ16x7hB26v9hzpA293Bz9iMnP5QOHq1JwnJbbhejw9iB4taSU+HSFsonHTzO+nhSr4ey7/eY
Ye5Sazt3Q2vVIrZgoOp+k8WlHz3RTHrt7mp2/VhOdDhSMoYbCiPT85fWtz3dFvi4Jc7odTwwh7vc
6NWbv/bIrOemyrOZHMni+uLvwC72FKSdDyijjCu/yOVqQbNWF58hbFs0hz783Uc8rf4fhzKHYsVV
V0L4VLhJrYJhkx8viavo1iiQ59Kv4mt4jWDJi5+W0Yo/yl1kWSROhR3DCViVzqZCeD+1qpJz4GzX
H8013Xnk0X0YcPfPNknWbBcgRCsUViCZf/snbx2nuj8yFm+TiljnZZxaq731tkVFrG+6mcQwpFLp
s6OJJEDxllmYEYiR/hhBVobaJ23hkjse3fHVHUNS7WvKH4ALGrVG4FVXvF9c8kO++qFj0PzJxwnM
BUfpHJqd5EWt21Z55v/F+dspb8wlC0R1KnBEf8h9gIaLzoNTwoxz6Hw35BQEZxLenvgSMgmJ8Koz
GTeydJvu8M2X1mBYl2em2cKGQEauAT05RB1kRquQzK+oWE5Ws6JL5Be0I5/MVUytkCkzmoFwXZJL
fjjhkoHSN7AgYG75HLwGO75cvzBcOIYtchI4VWL1PINDeyRfScP5LZg2RmQhyOcYj5gwXQDqFP1c
R0rMQ5IZWjf2JjqEm82ZGBOenpQma+4OOKOho089lRq7b2GUKEjiaiFJJ68H1FZG2d5j9msDlXSa
QDR/6NWLAPLLrrzF2xuea3DljWNJWUqY790gU6GHkw1G6HeV/xGLeEl3W4yuWO03JvVzcS/hQBs4
ReGbs30i5k8HifkY45bR7ixp29GO1JYN88YP7unp7N3eiOie7tJpMBlXG/MjQil5HfoLOtZZ6UgH
wblmFY1QfOEt2tc83Dd+yg442kuo6FVqxVpj53Qu+M1hlsgpmsPDU7BO+pA4ZsDApWoGbFLqNyTG
gj89YoaHf1Bvj49zPX6N2e4aKkc7CcJThFUABF0kAjQ0N/cKJCx2+k+eKK5LcsZADw0UyL6harVz
nb7k88v4cM/wB3wSRwPWHIdQEoaDFpUVnmNBGt5GBzMtUan0dbxRbD5TawN+/4nEjwbdutohkksm
2xNibC5qT93ZP8Ih0w0dN6nFw0rXAtWrF381+GaH5UYDZs8ZNE2C2s2QQ0lavQMhmOXG0qaDaGLQ
NhrLNeCDz8v9Y4z3hasLGmu88CEGmitIxBYwAgzbtRB127ZC7zp5NcLcvnS3uI4ebC1OBkbrkQDv
6eFNOYAw9vGYWrO8zsFDjt+yNPADdJ4d0EHmOQrOmj4Y4k239whaL9tbvjE12azQ7ymdJNqkdDCM
bcrZBza115xEb90NVxMWke/ATHedzx6DizgVh0vzmbC5UcQQYiZSYOtD2LONC2Bq4h2mM7eUS69s
wFFJeFcsqcDDeb/A8XTlmLonZfKbKquWxsHulO4QVb+JX4jR7eImJRyOwhRJvcos9arQe79s0hqm
Z/S6LZ/L3k7WIZISrC40rCLxbU5KVGsEIFXMRLFJEPeDDLDxMZ26bgIn22tbRKaREA4nIrHakaib
MV1YUUOqFmadBr0LcoJXdRmxGEZ364PecpWZGDBs6ez37uc//I5JYYcyguz3bjIaHaksXijtUEFi
aT7GKPNBatb56vHg0DlFmK3/VIjFunidgZ+Er/WNuzqhG660GpLQjPtrKEbSFUPymY1Xp3olq0ng
wg+0SA9LchkOOrPLkZEwl2KF2mAs9A/a2rETjNYkz2MV3HsQx5YSrT83ELCndS+E1AnkoxnJBIXG
YAP7+DLd0z4T4KRGoJccXxL//TiqONShbRP38CdgeNrujYmMWR+UVleQLDHqvfaUudMlMKRPBIfP
I+37gIHmnwy8V4ziMHEoK2esACyW7DzIOxyW7S8pkhSIbJDqbVORtkFKZV6Y/76h5VIYQoA7oRz9
zz+555arzEhL0nFKRGarywuS0djNvWwSbAKe3Z+AiomE9+TXV9IrKJs+n+Zpw2R2EW+B9mCdxcAz
1+6dKr0TOGh1BoSJgwxcWuiDeHzGN134105pbXylfGm5dsYLxB7MvrfSRY7sYdx4iUN9nwZx4xmg
Un6oHRepVvfGCIwaqC01c/NdNcyVOoiuGMMYKuRnTxW6CD1982Ufski7KPNzgXptw2dlI3DLBp1F
KFisiEOL/UFArVM7vlu3SIYT2tMLbYyQFh3bKJo0Cvn3+gxdyhI4H+lJFFakg9TsYkrmZmdIdgZV
fdZMQtB12aEJcYN5Vjdbj42XRr1l1LDa3mAxdVU6/WOCWg7SFMvvQlAp+xK7IOQau72MzAvA24n1
n6wYZJQHqqGvamD72VEMFY6MHSJHgD93CZcMf7x3vzIuFHDJOAvdN6xLrbgzae1JLJGcIKRft5g4
c4aPo6IO8fdvTxB0//p1g5r2J9aAUfdLC221Rb4lI7zRGvmpAuB2S/MmlgPA1t7OjOC+J7t25YNV
Yb/VYTFvcWVb9lUGyf/PKRa2CNQ8bjx1eWYGxXFjUzFvyPtsl56rfxnqJtI7iVLNBrvsOTsluQU6
bpuAVQq5Hzpd3ztT9L8oA89VSY8nZcC9mmXBlQzKhacbx1DvkxRi/JfP+PTDLoA3h/Rr5m1Apbah
0NEnt/A9BsXtehmd7DpAz3Eu3g5l4QbMWNqvGiXe/oxM3XWvU8uw+HmEtT4/JYGIw+mWMyc2lUM/
bZDIgcCCuJ0y7xi1mlvcPJOOkV8Q79ugX+F99NthgMorRu9y94B/ksLpHhQ6oDk0Vlfa6F8Yvi2Q
7BYKq9neQOx9RHncKCuzgUFIxiQmc9eA/NhRRNBJasv4sIdFyyVZDHEJTr3bSWjK2hhTkPk+nqGF
9J88xlbGlFkHQuvb540CqWxsuit0f3iLtW5RZQpj+DgmHn8Jbk4KLVn43cOnpIjyrg+3YYqkrCD8
C+U7WkqN/5pbGHXXmbrQf7GrF9Ftd6UKCbTNYiPfz8glpXZ2YXCdEPK9/b0S92fugFDSpkXluKqy
y5tjNetxj74N6E57hGzQ5Jd8YWnASXUuT8unw80yRPzK3EwMTUxG6sakuefxEyyGfwlSEPqDOdQO
N6rQPf+VvsLALwzuk1OykK/6KhK8RuN6+18x01iv1pnemSZN+enaNPoMNLItzibqVqVQNub1/ARr
kxUR5NzL3TeXgqRDJkuK5maxqcL8pyzCeUp5iLTOGzAOs1D1xQxrX6CnDd0VruEcHhYwWus4pe8q
rD9OePWzPm74t/ikEKzjGBkt7CYl8aD/HKRP9aSSd0tV5cMRtfyO5qK/rtDw3dpdu0O0cdB+d/fL
MJfi5HclT61PzAH8NRef0o9deYyxvE1+gt/NxTxnvmVKFjmZ+uoG7s9CU0veiID36n4gs8exCniu
G8xDNrECwvPuZZ74pFEdhL6yreMbN0QYNWGAomn6QseneCC/UkOVHo8INGWkMVuPNtj3h3xvrCds
PxX3O4VhuqEmFtbibcS6br3kO0ET85VtwvUMLBO1N8loxZMmptNt7zNOK+3OBgqaCRKadSkVTz+1
kt27ZidvJFmyRn5XRC9O3OdowpFxeE24nacdtqQq6+wL/g7qYTd151hf/HwV0OFTyYy/Ezx15bVZ
erZekn7qq8wD95M3bqYjEVOd48y4qBGav4m1uNAYZMSXRnnbkiy5YwpEJi5TeW/M2RfyifZMTOBx
A2DBKQzX75GPV3ThtbjWp8jk9DVDcow6BTZrMMir9fLqCp1ftVkFFAfk/EJG4IniFg75JP5SU3GE
RcWehc/34no/92tXQpZTzc1dNhnRKBv2whSgDpZriB3GfXwhprMkOxA/Uc3Xd/wocgTneUoJz4X6
L/HlE9kN3VWlFgdzR8RdVIAcuAidOGXcDZFfuW0p/n6aqzADxPauN/1Vu452qK4sokv5NAMZvfzt
hM+HmeN4UKlyRLSsIirThSPwrLa8g9y80MsqYNgP+a/KH4Qx0MCaDcy1TFRKektdYG/Qv6QPIBDD
N2/92YViQZ6G6v0lWuxPa+XGwzYQsLBhim2NEfBrAMPhcLM7YX8mNjdrqvjE54eXA48Q5v8HVVzF
6PIuIkE0dyrbjCzRMUiKihMuhj2fF4gME4FSKFd8tqvfGDtqbHLzRnrPdGGw0mJSF18IXG8G3SN/
ztkTzv7JwkdHUw4jYgsbNy5HVHnW+5GrtreW0cga8SRlicCmHabm53l3Zo/bQbBqt1ChfRrX+Zqy
4DM8bk9A/LfqE9EKwHNm5p6B3LinroJIPAcQSg20ggWabjOWvv/yLjiu8QTwjf+FGOdhSGixPXWx
jWxrHuK8/F5wBGiB+Lp0rucaBDwiAESTABjNmGGcX26nOPkSNgNaeICgTnQyBU6ufAgxxRTE18vD
2TR0Aao18Ku6CxtvMFKn/lUUXhtvv51UnrpspZOvdq0xsBnLCx6+tvm6gEGb+bJ5MgdaKEunFMfl
s/Htzu8RTWX3oad3zyDqT3U8iZDdLb15olIUxwZmOdXiU9TgNtr4aR9gQ+Yoc0NL0mM3TFq+kJh7
LZ7MeWE+3KR/1KTmQNUYB9CWtI0IbJq0f2HSlxrM/Abdpe2pfWhlaW6W7jqATvBqXzOxycFgOdPo
eEkuWznnfmT/OvbzEEtCG9rspSWvY7w7OuAQ6ywbSqx1yB+oFQX3aBTBqDQ/0N4pIvFCMYNYDqPi
9KsyW/SEbyzrFnZv5qJOhFReQ+i5jtfiN12LHbnbQBVCjBwOg9H7iohHZZrQb6SOGZW93eUlqyHX
pLvn2Oc7auvMCl4No+Zeu3VRV1BhgSTGBgf8F4Bj/zvbeKkuu0HHXiRVoqWupAIF4R5w9Q5tDscK
9a7xfXKYkbATfdMwYEFZcwHrEnr2axoaSgbx/PL+EgWyTHBCb6w6TrqHiSWyZST9hQGDEpCX2BFu
ch0k5Pfhhtu6I73XXFIuM4JirFTKAEPn8YG9Ki/GRwgc3y/zCukEQW049wO7OXip/E367xFnmZqL
cut0eVaOiTWPDC5SNzcIDmP+AlShX8J7OJrHeMYplBmNoRTqjzTtVxjB03NRvU+yQm44iIof1b5t
3AMnWY/dYqU9+xtvjvba2Jbrrh628PVDoMYZnD6j+5pcO1D4tJ3p5XDA2jPp4CQ8ER6HbQt1Ap3k
Dh5FnrkT4D5wxX6FtUbALAENC96E2+W+ARiScbH0IcKwTOEaP9Sv97gExE4uR5gU71B/dCRlyyTx
3kUtgEwyOKeVpcQPYqRx3tmBpQ6SJElop/8CbxheLz0+b3RekOyMChbyAjovI33IdMWgdPqsZZKA
hGs9KjOrCJPCWsB1nX5xiqoyLi10YGbd7AttjVTNaMRFCRucB4shxhOYwLuMjZWAL0+O9QTRRM7E
oq0ODRjAHCz0+/53U6AVwUgfBMW2NQOHQ5Pe3Ir7bZa34RtQP05NYeiwXkERC0uFtfeQgp90sFUC
c0lONq6bgh3ZDwff7uOzWmp3xT9bKRBqnN0lFIaRnC/R4zvR57fMik/dA6AHAeVB5RPRzgvXjRo9
FoXy5CfDzil7gv4brDUvzJZ56mywREUjiusOFZ4K0ba1MN+sL9SLL3dQoqk0fMHRC8x7WbnAEeUT
Dm3GHFEIDVggCboyMg3M+qH03OCS0Ygp11z9TKCIABJe7MOsith0EBqITk759qAddXt53DEU0Jpz
595Zd63ICFid0vsdtckOh31MmqnrcYRjFuzAc8WW5fBn/q7eOiFdJYqAEIkKLpm1sC/efTZWwpbL
o0J8sg23hUhupHroUmZP5tCnCMr3t5WF7HMrJlMY119fKJUzmjC3muJB/rAgn5WTMBrfSEkZwBLH
0o5m/LQUpoSe70/WoNOybkU+/fRieZohUjVY2uGLgRfZRbOJuxCWXDiCsYuHt2myVEsx/AYMuQme
m9vW3/2EWa4KoG6u5hvZe99ezq005cexCQGNqOn7d+aim8vmwSoPyY47FzAcGrpw9AnM3S0DqABv
uzjoyC5stWpFJGNXH2gRz9IylmfjljsrRn0e5i/kM0GxBmX5EBIa0RA8HqZ42FQ2ROe56AMnbTMc
BMX3YXxtBoWPBcgHSp2WCaf7+Xd71sx3H/5wUJWJi3n2xeW8RqfqUEEocQLtQbW3b7OAfLJ3pQQA
F/ypDIMRZjM4XoCaj/pOUlUn76UGJG4r8QoYSzGYCFc+aRYoaqo1Mqyj+i8TgdSO8YDE6NUkkBKo
jYmqtf7/r6UJ+yerOxItrzJ8B+T0O/73ZfOc6LydDtofS6MOA+zHfVfNZ0vc9yLMdyaZi+Z66xkK
MBQhKpQyXaHkUFo1rAolswCEpzO10SvDNfZdNNqbFPDB5IO5QlNQV6jwr5pnvkhB+t1jFYPt9W7l
/NSuHWBrB7hguC0l4TpzLkKJHdP6RvhkC545/dcvgqQfdq0IpBjaAeOkFA5XjL64X8MepGSeTt+r
ouElZ8lbfd/wzkFYwYAG0L1Ae9mqglGWB+lPp66CtcDzBxkIHWXnFstQEuGpXZfHAnrVf/WwRAMt
3yE9sGclfIgnu1v/HS02i4Udo2LzRik0sLmYWPGWaywfpXqdjWc15dCa9CYO9bCk9HtgNQBfdl/4
aiKgLP6zXpgYsMh2Dg+bxjkSF8xbLoyoG4wQXncilMWcNqZMFSJOqxD6/j1pLIL4WRRDk+YX+tRY
fCDwAA6qe73iNvZtGfnSPS5hXDpsY5e6UHKIoSc6L3/4KSMC7R2tGrCoAGHAnTZIv7I6pLWuIEWV
7yWbSHxQ2PnXEzAkaMTj4WzglzpBFz5OFuOVylgSjd9pHAzbhu2b+qrA7NbYvZCWHgR/Y8//Q0su
W2YDhXT4/JPQpVI//jppcEnIn+X9H11EzmBQgHIiQGAwXfIcw6vadt9OVgEwqlg+diPSrLh+ZSoK
PP17iEzqy5P0KrSz1NP/rHr3T2jEgqUcgXmbtcQP5TrvawvMJ5cAlUDCc5oOHtmZ5rbVVatUotSW
uieYYZeP7q16+irpE/oGTm44Mc5ObBYq3GUg5VBB0IDQQcOly2IQf3aPtcS29A8yWjFufnb3/OSC
Mw2k0ag1XoqT3jPmPoB45HPaVhXrnzVhq6c2qY3e0A0gzlynrnuMOqDkNet+eBNTj+yLyj1fzrnp
sKz81t0OrZCZdHR7gvdTS+h4aFarrUlqqJJLMkTmE+82ElgyrC9VlGgYIJbEbR6AOcteI7hx99vl
Ju8hgWzjBtaiZhwjUprME3vSIXDAFwQHOBFfUrg07eq+W2mnRZudMf0IYCEjy2nGo0ux3+KSehoQ
I/Qa3HLfuASAhz2e2nsgy2P0a0+7J8S6hiRCubqMhoFR9sYVtajIownmL3YjHOwBImy1lRdVYxkd
r+7AuuNoyF2mdAQ9uy7d2bgqaAzNC6Deht8ulCZjbmt5kEmEpMpHUVg5k89Zw5mGQTuy6Fbg/wFI
9Hic0+MI1NTwVgsOq/Y+2t902JS2kK5AvUPLf5prDlOgJgtPs6oD5qllwAnUkZTfZbc/wP/10CST
g++00P/QaoAOyCMrJCSgK5oisDHtQ20MBDINgqTdV8Sce8PbfeUfhjmZlBcBdS6pNiAMHfaiWKVM
UAJsnG8CFvOK+FdR1+JC0knYCEAFf+TnVoyQXHVtN/5du64k19dhCpeakHIhB5kiEMMVzhxYDYI1
ckgLAehvy7wdYtedG7bKzIfN4lFCFtRH069AQVqdz7qLrG5bQo4CQw0D00KA/tB3/r/eCVBzhR00
N/wD3QqW5+EZVN2Q6s59UMXqrqRUC02I32IPXUztgnpH8f83bgcD05vJ8ESuAy1VnAStzuoaiyFr
mS+RHsWWKSTCUdpNn/ZPDAnFR8+J3K4yb1KYwEC95/g5sk8BO76OQMaKokwI78JfOkpDEa7AjAV8
zNcZ0N4wbhESsRU//YyN4JyzUqHmKMb/GLAVf7CSM1ejgimPSmFj6AIgkR9zYwR7LLlYVBBv/xDt
lT1LWPWBo3kU4paJxKPqcQTeB3/ZjO2AVEjFvpVEjSKKdluBmOwC5wHkHaG1t8qcZw9rPdgLsvo+
DF/6L2s4yaeEcj6Zp0dVkliSYZLpZo5RElC3Z6m0XXvc8k8uJqx9LR0uNxhY5jNtJGL2A+wTByMC
Yvf7iRDPZ36b/TdW/WL43k6eOAEF+ZP/KL7ie3i4geGJUmrw/5plsIb3QX00eJod1fatM9VZDGxt
URVLwF7+w2zN/PvZrtwNiCT7bDdUlocdDce6eXjoSyZ3VE80KeppQMAH6GU9m97ta1emLaW3Cx73
QEG/cvoVdKXhEBmiiziYkCLxfGSizQEMdXsX0Hdgli2USNF6EA06Gp3TmJ5Wtp9Q1R5Tuhzy/DMz
VMpr4PecMlFeHbiFrTN1aA24bxfV/EQb+Nw4gUAGHlHnhRVJLcL6dzshpeFWiHI+s1dkG7UwJrat
EcuSO1JENbQWpCOG563o+hbAcmcn/nxwHtt9pW+QukOwclJJt483ZR08fbUwCve93iGxrU/xoQbj
6K5o78KjTQVcCC7xhK+AclGrMWNi2v10AX/UvyIdaNPA3mySZ8f7vErTZ9CUWXpglOht02yqEecH
6Y5y2WwI3/LwHPrHfiPyPTx5yHdhjcub90XsQStC/s+0i3JnVSJknNSLbh92CkVTz/BJenCoh5Rp
Ef16xc5w4dvRpDI4Vvs17m7LgFUAFdoV7XVYKl7gk0lIrkGZO4zmrxGpWHtFGo0nE7WvB6joKKhF
L//EYXeh+Z+zIy+bbbn9nWPh5MkkuCybQZoPek2lF1OXtq0+WW+Xyf8E/ai/R/uGxMAmmkPzr9WW
MAEFCALviFoLJoj9ZebKYWIJa/KnFO/krin8XrjvcngEY85fnsHaQOSvYvMWgj3p8evL4pP4HawX
C3s95RBWkE5DAlI2qlVV9dbhfmjTOAa4kCTO0ygkaQ+EVhBiTRil/8aHeSKFko9XgADOazDvpjI6
AmSVx8zqR4W94MvZS+TeoiSNy2c1FgHI59xLmRe+dmkfWiXX4CV15lPruJCp89MIBYfZbpQikvEC
fp8IVlXUniskDhcMKCPtdNLrB6iYM5iHiwIKShQEGgWXtrXhPx8I6Gw7vd1TNUcDGsqjESSIb8H7
kvyiqB3xEIdBPBLvQ1d7mSxI+KUx3ky2wySflLfCeERi939lGlnG8tgrUjgS70FDI7ufwoUzb5nq
fuXMpoUNbsn5JaExKrihX9eLwFijGUWcsy87ZLPkjVi1PYbZKj0yELjEgPlGumhtOb4xDtFDr9w0
e3qK9z6UPh9uJGQ3cXLAzYd80zu0qXOFRvB8hIIbnrG1kyZ3MM5XUy6C9pbRCVXUpKCTItjptb4P
S8mziV/5rOPruuYMFZq/ayblpIgOa8RDFYJMiHu+heuMtfcXNNY4Q4660v6QWDS8GO0aMrk/uik9
c+TImbYDFlntufakZs1rom1d5cywzsjQEWvD3OWFkAtFYb2pgrSt/1sFGrWSyrZbYkNQJFLO5kJ6
QHZjOrgDobdYN5yv4ggmXYjeU1kqHoVSN2xQ+lMf2UekYsnfSVt8LAbkoL1S+pyIxZhnS8faKtWH
zTGbfSJJmPghM8wP8tiq4+lFBtdzBlexFd6AOM5BG7Qabh19h/t/182D9ciEYhltce0Bw3cG93rQ
LlNJI1J4Y1ESNQwawSZcgmNytdmtSM//mgRHBmoBb/0Jnr3n9SOMv8XE7UXd6/Fko7FUBUoXpUNv
eJZKFZXcrDtq83KMi09yP7o7Q0lA07ITsGHB8P5P/ryL1IhBsO736iUFQJRcxF6XGmiNIY8ZTX74
6FXvEy0cN2e2rOJrMJItD0StPsT5It3T7uM092UZ7+TLihq1EMfUNTtMRDPpxBUxW1fVEaHUqMmQ
UfYjtZgcpQoSxRikN/FtThdcre+JeXJw1Gyn2zH/P5HtO6brP1J6a/bML8EKQAwmBIRaJK/8R9AI
eEUfRqcbRc3g7bYY0J2rBGkVy6XvysXuF5TZyNFbRUF/aSaxyDgPXFyY3hIIV149l3I4Z3Qj/nEx
uF4kmVB8yB7jY/5BNnxhME6YpTEpQTOAyzCELQJo5LPkUGIYHdDl2kmyTZUO/EYTOC9bnUSNmFCr
yLxHj6f8R2DXQeASMiZHMycDKOi6j59xFhkfU9W3Hr6+ERdeDM8+FmeY2lWe/AYrv7Tp9ahf/VlD
f3ZXJi07oGAnTXmRi1JOMcqW/K3Oo88yKwKIVXg8miYuQb0ViCOGcPg4h/kVhaN1veQ2joAKvX8m
In9711ZM4nmO51FJe3d18p1WHH+vyN3M+1SA7AAXgBoS1t+1IFuLn7S6Tt4grSvqW9j0+tRjwhNX
tNBbOisY35pAEdyoEGI9k/YejYzwXFfpXSCgrStUS4UdIF2LpUhBy/7Am3IP9hCkO1415twdRMAT
pbuL8ABPiuUscYC5/oPC9pBMtsrRH1kQOaMpWcb1oy024aApOKPjzpXogbqT1x2yDudQ2q+5I6Cp
gHKj92BmTrbCH/ZwZ+WblR8E6R10S5xJ+WL6dYZkR2kcZQxnk2NdujBoGDq7FR+bR/7u15qTqqQj
EhpvDLAr4CmY/Zw0ioxcOcBwh8Z2IAd2Oe9Wl1hGvbGSci7ElIheoVvwoJpuY4zO/EvvX/flN9rB
KiDT7XqYXbcXCYzUUDNSPbWIKp2gHoLcZi0eMHtDNBnqWH12OWPDzA7cmPM9HH3JgWX3smfxFaFo
+SPVDdT4zt8OAK3IqBgfRTIUL57s75uJztZlXzMGEq1MQHtgbDvxS+dT294DIDHBlQqs24yet77m
jGDetsZQq91dRca2zsrqiBRhFQIB0I2Shs7G0+2zNWOHGttNIHSEj93nAxiWTPiuOKe3kII8D+Ja
8kABqAGGhiS5Y7osRPvSaa59Xc66T2F+kdi46+FifcXek/Z/U3gFyV+H+KcwGb5ydBJ8tLT43FGY
4SNF9CwoeNdvp9KCGkn8PxabPgkBp97+mk5JrfZpNFV9GGZekZGfxZVe8fEU6a4R85+McyfjFh4P
abFdljZ5PwEW3JvBnRPW5AmkqhqLPGBNTXHmIWpRzb5K5rVz8jz0pK91YbH9yfA8Bw7SMmUei7V1
2IG5PLmjqtSimX2575wXonzbdlHNGWTX81XnU2ajEU5u+fN7vfvMKwCfYS2j68/37JK/p0Hyy+yc
6OGXKbZGXktedk4kSPkhBJmZOnyD7jz38HGMbsCSY4bt4jwxO+jJ2QWJGDSWrUcu2c84ARWz65CY
XBwaYOA5XeFGpVm5vAExR6zMr/9FQ/sYFYpmLAe+9O7bQBkTr+tzp1aHa+3FFMaT9z0PaqDa6eoA
9BQoqW8ktdgZxjNAFGlUZtpRYXFEgMmYqCMp3h5ElmPPe7+YyftKe+vdCbH0tQq1M1GvCSfVX5Vu
OcSEkyfzPtuj/bxbLswKn2t6RguVMweUoodM9nUNcPKEsee01ufUv0mGXOaqFhgb81gtbwb8n2+X
CWeR469Mux4ZuHQAgYrMf/MRWXrdiQZG75eHqSFOx1lNk6SqeCZ073QW9iDk6omTmsyKwoZXIjGx
3T2wdeMA8OGx11QDRRu5rxtt7fLinKwOXZUMmPp+H0e/izJp3sEfnVuli8XgwIXIHpv7j5NFiFAR
ZOvbeO2zqvYEeE9B5hkvv6qypFDGxBQjFEbq/U9IbymI6wZNzR0BmAZlisY+VAIYhGuEuS8h3VYz
tv7tihCSKZzDHFLQHlp9kByHEenRC0zqdY3J0NWr2n0oS7Y7suXvxv6FCLc4EGZhXycWoKm9Hi3G
wS2doATDAGMlvOn/4RdiEzWOCsA4lOkkP+6I6rhgdyGo9RX+p4yM6YeMQa7GUocPAi69GnXgcjkd
FDndLrbT3TVQUsNGvZXA/aegQRGTOS9/guImqIXU5vza52rMbuZhgJelZytCFBFRmNxQ97KYTyhz
Q6inF0WG9zHf55zn4fikz0V0/D/D3aOLFoNUKLehWl9UDhutPahJbpVuSrpzZ0wfLI9hhPT3Oz7N
fqXEuFf164v3LS/fAqvydagtSM5o6xYnfuJxoRYXl+BozMQi8R+0/WRIS4/DYNfeM890uNTaZkXc
2p5yhq5zX8bBSs5HSOkG8Y1dF8fRHJVgvqpeBewNiKCGrMiRcVlNTucznGASKXgbYXGBwQi9NPFf
m+lVOTuVTciKoXNXwAZ70UU7xxDCn66+lSPNJeb5wYvQPr2cwuwjq3xeM9vRNn6Ck5Y1Z2Tyz/HY
ayj3/V/ozA2iariVXBng2VmYlu3ioL9vS+SWMgrDpM4Riim/dY2oXKUuGlec8Avhu8bSbeyBDqAJ
aYSw5RVS/JbWcPeEfEV1O5UamwhHBacrdm8wObqK1LR3DbD5pQYyHMrn8ETAbX9t+QB0xv47YxOS
cG3YZ1zXAbfrrqsFRQv4l7WciPhIEjikcIzQ/iYqqAcKKn43sqdFtJ4CWo1MrWfVrq/DAAfRFrfV
cuYk2SYMjhcvYK2OqP/YDRyMfrPVUDsR7e/pNs2G5vI7xHQJ77JwKTFKIOeknuxvSTqGm0x1p/Sb
df7d36e7LL/Taw63gFbv3I/p0nYmMhj6+JRrOXW2Sj9K6bg5khlii4Ehz/vpUPE6ESFsvySnG3id
WneLnIibM6lBPpvIhf8PrRDpkChy3BeHRdmDX2HlzzvUhe5T2fhSvJcXRmnz4mmYMXMjDQfuLSFM
+nrakXxJw8nMSy2lIvF2dQV2ye69Jl3dcsaGC6mfhWQ3ypYh6pWAqWWe+0yB+FoAwEUCfpjHsEKh
Cw4IM8iM22dLS8i9v7+H1v8IJGiPjOmmSq8O1lHnViGenL/MlMXT0C07naLQXKGvZKZbMTN5tnrj
RZ1p+y0zzn+C2OpnhWsts2E1qmoETVvHTNwKN2mObcsJxbvHM/BFw0UYZlczVpUO3ohezgfetRIV
JSCBsOokXUKnA7sJ6ywrlRy+lCtje36JBNVB8hBaUaDqenBRsM4Rmhh2+NuTgy855fC0lhZDsK+A
DUI5FBcYBeJqF0XzgF+iwg+Xzd7p5Sc2SjuaChcBDtj8UpBl+TFNsb1B0VNgpKGKfWUaBdGNexMo
hrLkDP37IyIZQsV7LQoVTUJywjvWTKxAOfwTloFBNVESpZvmL84CqcrZN/l9Jy4yXizh2uPiiE9h
da/3T43EUseCDYIizdffGa4XG+g6RWF4TRgIarKs+lBIgulHMNUv/yD8/kCGVnbD/Fj1ckr58ESr
FTH2km8QoAi2sn61zAIQhRHRoiyx7XqXW5zgGIr2Tv439eJ2BfF03RirQiVbUSR/kCaCtlyOmGNz
m/TGsHw+riR+dsJRqiNUv1A1XkNy47LJFSXiS6YXmUIAwkGeLS0rcirRNIHKaOWx5lcfrmP4STnR
hRQxTxUOFI/07wdAqzjEzeT76aViOIn45o4JiaA6VXB5kCiDm4q9jIvnUYpSKLIeCZw2IvaiAy1/
TnjuknJL3nj64P5uOEnAtGjkvoEUVrbo8gAKR243xZyHcSbFPMl+XOsz3Ou2yANB2TWY2QoijRen
7Wnbnrb+Xc55iIfz7QeMBFPmhTV4R4nauWBYW42QDQzNy9mROgfamdX2z/NdfZMXL9rNP4FXgWW6
cHU27XMOQW4N6zeeZNQ1z2AAnToyKzGSlCfPAqRcD1Ac99SaOEd33psSVLZL85emeEp67GnSolWD
jegHkkjzc3TA16iY0iH8P5GY/Wh8OMnSy/3hoF50qxBFM3q6fyiYNqIkHkHIfM3QC8Fq9pv6X7Kx
iJ83Hy5ifT3Jey2qj9dmlXa8KDQP0bpiiqhOVeerJMOvLbUoeDL7Ane+M/kqsLtz/u0fOscaAn1V
i4NtGhXaQ2itzh5eqNgjfikvaYID9U9G4Nth6jqPxQzAVBs21iHF6yu5fM2l8yTIUn8Zb7/2thsj
SiSpQxvM7cUWlg5GI3sRCiVGlpS14DNgX/fyojkrcfFfBiy509jIm2A3JaBJeSd26p9Q1Hn1q6o+
QDuCSCNiAAv1/JtxqwSaUH5l3I4SsIbhhHWj9D34eMjbP5NfpnA1a69bA/q0BcESN/6+EINT2d3C
gXq9/Ttj4WgkYsDEP7A0T78qmDoBdfOdvvhuo8JOmzEe9hBAiN9rv5tYHYfZl7GIm+oPtrjHxZVt
/CAFEbBdXk6MpZ8IumDW/33ZGdZGkcNZLqEiexh6gxiSOlja/6Mn3i2/1c9ZfDxVfxi+N5Ne0dd8
JkdMP+V2kf66hqwWnLwSECL67D/LRKVCTG30xAAg5kSMlUYgO05lOmv1VWWrfg124FozX0IueAGJ
AhalZMPdMn67ZxdCdUIT2LyGuocujXRWeLJSGfF0Z8F0c9BM5ABrZgzqU2E5Ab1v0bEhsZf2Z89K
ID23iEnIK9dgACZ5EJnxBwVtTl91SHfEqoi31rp2TB3zfK+M60eccC6xK6lWjdvsMpD+iAbGAxuP
1Q1cFCt1UvTLA543R0nU5/5sloo2A/k6CMqqpBH+P1erYO9fhB9hVtjKji5A1gkyniY8KCpLmNf4
ClZ35q/8AK/sIMJA6EDVrouVDyxE2akqOLRLCM+Lw5tlp/cn7HXi48Z4LUI3v/EPJRrac7WnAlQ4
fIx+gmna419pqcXsZuJuFVu/xoTGe3SsJC9AAQjIg5EEmk7mcjBGGRCi/LODUu6Gp0u6OxLQPHfx
t5JyKhvEKk9rN5xRmU0Tq34SeHqcX11ClXvJFhwpaTKTje+8i+C4sCMo6fBojd2A8Zm8zrXzq8KL
QgJU9fwIyJd2MVAR+QCD053QEe3PvINQaQyBa/RCgp2ayPqYVNXYRAsen+IZfqYvUnTQpWTb1/G7
/3EHnYSNnf6i6k19gVyd6b2l73UnCkX1Wi0xGJ4Sr5H0whCXH4dsTPpEdcYhb72nmnj8A07pLVaL
c+15hfkueeSy26aCrk0h+rgQ8pEspbfEtFIerD4mLrE1OZkQIqCsSMWmIoXuiUYJlZ/Yi/l6dLe2
P3/EWsjUXFEHlvybZiZd8UKQjbU9w5HEoXz8GZoGiVhSlyXV6ydCZH4jq9tEqkBmXTC9rNesf1eD
y6E5i8d39AKPpDkCIYyM+9YxiAdDrA5e1EcuDbJcaYQTXEI7PBGePUzQxk3UhCJUO2KDuS9qWpWS
NePDWw63H2UvykyUgFtaeoTCRiLh6TXfYEA+lDIvPozdFojCDGRjq0U3saSZIB6+fezVhXL1pEH1
9WpoXHItHRu1clW7/4k7OG1wyyOgYbtG65pI91lz2spr6+0n9IJBMwVipsU3d71armuGRikOqQum
ZmWCPyJMSkjNjnPrBuJkLJ/J4J4jZLEobynRDU0+5vhxxVNux+rOVU+1CoABVqPjFjG30K8e4E0K
j7fCgCpSohD35Hn3r2RHA5VSnXofmYTPXVIzdkSQ9mRVW5dtK0VxVFxf5Os8rplyUdHFqCsvD+GK
QrQwJSIfpsRqAH04ekvUN02rh7Qhw75alLH2AzjExRKFmgomaaCyUV0F55v5vaZG7Uf6oKZRcAXi
UoBLmNMwGd2eUQa1vQ5vQgzAPPQ9DvZe/ciYi6hztxXsVPj2zwRHqK1v+yQ0Z8klrRBSR2GI5XAF
WjA/+edeSsl88ZBnCIgsEPGLWzYTiD26rHPVbAmAdTLemWCdzAHC1K2nhdkwkmB/9IX2Ww0m6QFi
bZfQ9YVhd7R+cqr6RZGYwukDwdaRcSZEMXlf136LTr2Ml6YmtIaujOZhfH2chdXC/S0mBY783Lnb
otLkC85VGX+0JWApkLHwiIjDOKSj2Jh0ORzDQMNRcXEAeIfrjjKEKbTBYfyFmBKh3iXZNP3yR1eD
7/NIaNqvq+OV+6IPvdSqQytzcIySKXwQXGPHLuxuhyeXJ422JMSK1i2EEzJQwzJiQSKMbAvGVKsO
RgwMlf+nZyfz0bkz3tzQFKmnZh9M0U1bOEQoo3hkPBeCo0UPaLTSNYyNNXtU+dnvtZdu9iASpkuG
xwli/KOu5E+6WvnxFvmuRYknPm08GfYhnTF0rDvB3sILphKcvhmNixmEX7olmX9+gc8vVXLLGQJf
5Zl5r6BLkh2UJXEpZQptTUiaM4s3aNeTJNX2oKjKHy1fOhVWP6UkVYSYo2j98BfUly9AiRsh+xQE
Bj3LiA58FTBUvBjCi6vhWlPuoNmdtfemQ/FtBes/ONsnb8Pk3qTQOoiLl21W9U2VJfij79wd09so
ZMfe5fGUVy0OV1jj7/OPmxnGzySEzBE1ciK5TQJSNn948yVZ4iIbr/o6S92YOUQRXpKzdSzyVKYz
yquIZaHuamaJ9uQZQnd2Bsx7LwPOY5WC1EDs7Vb9gmmprT1DZMKZQKBIYLJw/7jV/40G8e2xIj9e
MtoVDi54A/p68hCCjvJhzcE25sXhmIxcqb6enr9FOJFK+sbB1iMqELSeA0F//aIq0/eDARDTTdGt
HjdNDkRM0+ZYf7WX5XkSO26Wae+r9/4h2suJ/SPjf0YOheIxn5y5Gm3qgBnPL/e/gqDOJKfr3VM8
eWhquhVNd8FU84btYwmMto9owDXJFucdjw+orTi56hkUNWGEOeAegq4thQYvAZNgUNYEoHjhbRlx
MvCZYpt9sf4YYHsx4TAHE+z3mBuP/iJHE7s0PKev34nk9drInoQb3zbskYjcbiHLXf5q1GJorAtp
Z5MqBUYHAuVW9sUti08TvKrXIJrVRxyLSJye9MbBeNq4PvECc7y55LDSzgkuta2d1eXo0aDnl9Ro
BEV8tuvZqyiiHlV2WQfNQVID1fSohDS/sOgdtUlbKnCZ+ysyMgNVOkTTjhT9vJ9+U8lJzOvgfSts
GrRC5tL+TbxZfgMxzmkvpp1X4shyNrT+IJafObJ2hraPhITYDeDJSnmGC3hHsEaBQi44qdf9CzZD
XBysMjbi8Sgh4yv5tjnDBip6dTzh3dCmySOfv7hh1br7ulEMNMaWoPpiDquhnGkkKKWMkBkX8aSP
9X6GdA6jwAnXRly4wrK9buWvbK0W8htfl0+sC/2wbZKTr1AcSWp5ZAXMY1zuE0GAKzNc/BOp6/Cs
UiOZOFAf9ttWUNTMD5uOPY1z90x71QaTiyUp/qM77enEwmJekqq9qheqMiRDO0qUGMOYJqictq+p
nJALFVAfI+PoYCkfWpVTNsFc5UPagiasCsmaQvjWdTV29lXl1LBSHB7YuH+gT+t54gdjEuViszHS
OtBwDMEDwk4mxQ2xst0gStJHdt5bvwKSSIbZU2zwpFPgnDOdDNDav2l5T8M7yY5HoLOPCaVYNmYZ
4EWzhOlSghiPslVcEYbh9PCPi2IOSliWGPK8JYKWwh9EsVAp8NWx0vw6h+8FDqXIuss9wVLzGKfb
JCQ0MH6v6Gmpg92KcRlE7fiYzWigFzmgo9c793RIJcDq59RsJhWo0zWgkZSWINfNSvnaK8nw6AYg
J4YraexYqe5cUGprGBV0Bi9goR4w0pOLeIf5UNNY+rQUuMVcJw+tu2h/v6uaaBzMTQWPwVdF7t+7
QFibIn7WDkuNY55UCZwcEorLYAq8ci1w5zCmT3biV/Jy87mC0yKNq6zTfLnps1n057YpL4zoBQ5W
ye0vh2gem970PhnVsQNpqTKAaZtAyrbr+FXNd/oMcWCAYlXXQR3Q+pljssBjcN3gYEpUqtjAYYHm
pZlsaemBytS1dnmMOR2RvVSmYMZGzvsZRakORuNQeyJpAVx26Q+DIgFp5CkZLfyOEPuOW1cIcqwu
W/i9EJnhale0CGJ3Bnqq1YyorvVVcZiB3Ok51S02jxb+HPPRlymY/qd9mapS+RJsq6+ErxSiqNhI
QncFIxpaDyqcTdiAUPecdfnn6P/2a5MzRgfJrinCKD0c+TUbVGAmc9Uxkit1d62HnlqKoQkALRiA
1Si67YkYHdMN4kywqwQsTz13EDewqEwOb6LJmNqHHMuzpJkahJ/PlCZFeCoWcKcvBKHBqgBRplBV
BqQn5kbQarFFg17GB77J0rmTklH7fWpsH+dlnkhmbopNDrD2HqmBCmNTAhf23kCzFsenecH+pIb7
UkKEipXbH2tZ8vcc0m4vLd5COpavu90Te+THooSzH3vXBYu9Y2442TmXpO3nY9qhfZk3FV6WtvXQ
Zs5pMtYf9yrUGC1rZt+pswDcWmZ7ebpwrVIYmOMaXw79qIjo2UFpvsAQbpaSgsGcHsJCWGiOh8m9
bnnTWLIq09TNEYLWp0CyynjwPvKmKiKqmFycs17Q8D++n6hZ6G1MF+6yvdNz6yABstuBlyHQmC0+
hcPOiJdQHtHpw3tm3OTPpRGLXqV4Pql/02fIP5LYtkZe9LuUuFX0d54FO+lvCWm1Q1B32zCCrFev
vcqlNXwsw/wRtc8O9sKOS2M/BfIvBRcPz3Ea7nNQutYiuMmWeP7WIeIYtw2uObk1Otg53g2esguq
hqvrDScoeZDm39bBgtKhyvws9zYdMfVK+KeOjj1qfQ+oytf86iav112TMtJ1TpmU8w5TgM7PiuKh
JlZ6/KotmK0s40bAB2OLoE2AD85xf1wH6i0vGGZSZQYu3ME18Csz8UagflNDTB37/CuEFVGbpgoC
PfPE5X0ioFBwGro+MVHfYbyT5EWgyyoxleOtyNPgEd0ZkloDfgW5/PeQy9DRl5ZCmq9roGw2lsxU
fddw7HefHD2Hg/9BWSZPqxh2aa7xmAPGYyM85//N0WwtGaYGvKmjcgVxOnWMT03m2oGEX0c6QYqc
plhMxCPuuWKj3lUhLaBEw10UnO0QmNpOAoVNnBa2PCdtssLE5DK2DYZW/2zdKTG5Drm03w2r6gr1
3Yfiqxk1pcxWo0l0kNnMplYnwA+vvMwyWsDU8Q2tVTRMfamch7wusr/lTLGZjnYBZObL+BF8/LTr
jmAAfFHTAZjSXu5HANavBrpIg/fFllD5DotEja1HIHfeuA5jkj3DtT/U4LW6RQRkyrWB17qY4YM6
kaEYNk+tNgnS0AxIAYQlN6S6peU05zbPRmKed3JcxdCnhM8q8kiUktTOA5TtuFbBzs35dOxZghfe
4Fz/1+C4h+WXGSoQ2zQz1leg0bks9bw4nA80KrAAfPcHzvOIWwVkqaM5WQ5uMrMHoBIuricxHm3w
0VF1Xrh2Z1xeYtkKEkyy/hqZQiYWml9g3VeuQPLr8JP9ImoX+30EQ2Nq3ycRclgEEWyMmyBnwfqF
ygY8osvipxIdc2g5e0yvt1Npgrll8XWOm+/gaQ2ZZAc7pQ4Zu8PDXGE/MxIt76JoE/iYkL70EgFv
2tpmkbK3vR2U0B0cAqZmXt4PcQTQhnFtUoQ0Dr+f1kYJp7E74K8H1jRHh8ohuNpDnj5uAci5KZtl
ImQF8bwKJKU2i2MlJTv0CqKqJqjnJMwSa7X0ySQpzo+82P1L0YZrXHQUENlZH2Yr2L+EeP1FREO3
n8sTN33og8+eeeV5DdZXK4A8EkU8+PYSPC/Ruh67PfAtVc1fJ4HdZST44L23dUS2xaC0txpTZDav
UoSEwWiv8nQpoZzPr4fE1o+ljHeTEd6XRVvo26NA49nnbSKK9tSMTeezcs/aYGPQ+BueT27auUN6
En3Dynb7dY19nWVXtsAV0DUDVWKExtzve5NcepNXTSdujBSIFX+DlLNKFNG08L/bghiR8ywvHUip
++v+D3fwKm0sLUli4NIxUU9kcVbTvklMC6ySGFe8P1O1G0nHx2YfQU11hklZvcBl0sdXb46MJcVO
8Q9RlspvOSHm8OmtMQ022MnZciPnzVezfeIWiIRZ1mcXXAT+xfyPb02wTimR+IUC7JC9aMscvSwg
HlMCYOGGWE5PT47CO+6+oXegD+K7anL3cFe1fr78yYQx/Wi/K/TUMEh62hgJtaEkuRXjF9K9jtjO
INx3cjwxQbIyAtqRpSoATPlxDZkrUH0yhwqSCQZFBWOs/yrn0OonULQ87CYwOFLExh7lVrpXs7zB
hfO1aH4Q5SZwDtHbH3/FJGIcOOU4AX8IZGLDCCQ4vVAOqI8w5PXoNdulea3cHzy417ho9pNwXBS8
MHMSXYX3C75s6wrcN5rgPhGtocNppQ95i1xCvWev/vAh7y2pE5iOnRLealeBV/a/9zQbtwNaKSjo
F1sDlWV3zYykLEQUkzaS2zjv02764uOl8+2qDP5/Oqw9yJJpLOp+Q7JQBe72BMPnE/yvtvvTL5Q/
rTnTQLcKxBxV7+5ZBASCb+jdCPgzyPYVhPpauR6zFlqLPgH0IQ2Xt9yR+8ahaoElVDfTtqlkOvaP
1WEs+RJpo04bccoyP78Sck3XE4anu7n76zxu3UXTqdwWdzmjB7XMWr0qiDTWZbbzgiARvEtt9p8k
3aArRbWPqfTIon8EScWzqqSuaX0eLk2ZlviCXrkGjt2R5tpseUXWcDh0Z0pMlojO3OtHdXA3W+Va
Kp/lOvwsdsU+kCg3POl6KygxXogzAbAWnmTOjrL2shpNeJIvb+AY9zkILGAOl4l6QqlQ6OZBqovC
t97EX6Xc09H0vT35yQH9WZQxZ6sQ8tCQ4PNlwCgzKQsZctWxVJLIl5ybdgGIRUnizAiGbGEc41D9
K4tGteoeguYm9/hoiFBRkOTQkl/vfQz2ZH1j0gKCPofE8G3JOU3zZui5NCP6gmmbSQMJodSZ+ZlJ
7scLeMdGU/AOEDjYNhNhRcagIiJfaVPcKJt69/NRFQdFYhqYgyhcIkbSYhJJFfkvooO1aj2Dwpw6
soHoIkG6NQrytVdWpqznDmzXYgJhpDcnJAACAM3MEFgMU6x/7+Y8tf0ptKWWkS+SN+nDo1m35XoE
ppAKNpEs4mAof0bXChmKOS6AaUgBTAhPWRhjkuPXiHcQ6WMAcSkq3eCUQcFV1jrHxnH09UgZuwIV
OtH6EBAc5kEAIAD3+sKUvZ1FR3jgjnjLxmtb5hnAtyTgAXFiWjhhEo/LLnQHUh5LDykE5Veser8T
K1Td0UhO8XDy0XLbJisSs6DaTkk+zJ5gQZXlKoE3HNOp8koREmgJ9mpCc+dHQ0nBVfBIzHz+lIu5
NJVH/7AUuy6iJtUwdka241F+GNsfhOvP0LbAb0dQB9kyBepYp3hQJJ7i9Ux3kVLX1dAVw/6uEZpL
AaYnyJB9XyBQK6cTZmvbKb1sz/ROaS5KAQmIuM7wg5dBbew7nwbaYxneRsWNJ0VkdWdOFwUKBpb1
wba9ZoWnBCQ6jDZiUFB+spXeeXn4u4IGBBKeMGI38AeFqNCqUH5iayJ6gAesQvEhvLpqi6+D2swv
oiNZMaJkJgxNB3KUVkuVxRX68GGIU/A4mf8PE9dlcYF3oQ4Jl635RdqArCvlBGXdZv5KwqiExj5X
O/suTL/GWn+/3rnPlZM9OLtMXO1lFGuyD7un4htoy6izhInwp+DgZWAd9bHzzVEAZntTxoSNtuO0
dBAPjc+YwcCk5tCzdTmg0BS7ndvc8z6/5dMDhWDJK8y8HRuaBbX9vz6+odslPbektvEhDPwesjjh
EcCd3GvVD/FMAP1GfvBJ4EBwEjhJgx5i3fodns05+gyoJvqprrx96oVUK/Q4o/1zw9kHRJAGsoC3
e5oe5XLNdmmyou0xQCZ7g7yOqTTboHWzTu9kem5CgJGfgS9BWFqSgVDLhvOJtrk1ytFxq/E4eZvD
gCTmMw9YWPEw7UxuA2aXpB3RDWpRAtGYClRG4G2gpPuwawbG1NKtLiebvEX+M3UF94iMC40JSYR0
O83b/rL1kaB6eQza+T6iIBMHNuE9D2RO87Ts1yVmRwKB15Qa06jI43fl3nIAloKS/6BoZ8NwR92x
vpAd2aSgSm35gTP303DzNp3lTHvyA7qeL3RwZwpLLPRCVD0A6wkmbsNkxqKWy1fb7vZYOi7gryNj
2UbubSLu33ivUDpMIwCBfgkP1cRmUxxd2ZLFhbgiGPkLZ5XvpA0h/NqoHcijYzxDdHkz8hE26j66
ctoe9NXDeVPPOKwfBJZnOExZWpMUwE695vPi2fTKyrySXrd9fgjJ9f4fJAFlpm/nNDyLkMpXlnVV
pOTEn/JUrtTUo8K/vqmf5k3GynWIsqDcdD3pHL7e1BT8MxA1BIPANRrAL79YeY1yE/wH+DjbEoef
moYDnNWd9XQj0Lo4kiA91A0QywUs2v6isxWr6cjuZ6GYSP7ppyBVQD1x403W2mDWuPa0USaL1s95
Ew8lioV+kF3FzcCHUPs5oUX0nJaB9YIc43sxesE01lCXPotQdlyeYkvqmuKl+KkDVWsq2wLO3UVe
aBxWEvzEdsfDzcDiCSkTRPQpnQwzIH+lgDtMbFSAfQBhn6lEm+o961oZPUJ9tSiJGBRUFQCEBSef
s0g3FUflj0ZU/HQ79JkxJJWyo6bTvIxwjuqlaOUZF7YQkcIyOBRTG/BNZbjvXwiWg1bztL+Gy/WR
O/MyH6kZQyGj2R7EvglPsufGsUUHfhfA5ekfyCXjbGDH0j2betqqxbAXEJxvyhIBYaCw0arhx5Pp
wuW8PsHdSISTlSE5y8tEc69yrUS8JIGFNIA/FeyD5xYf0DnsQELQ8yc6EinoUydE0i5pfGbXMJ5U
odWd/5pjBjnDlWUKE8dBynR+m0xCwf8i2uU8jWBQzhmQMz9Veg8BkxDksD/CpcuuTIGy5e0ECKNX
wpHXsTdqA0VykxQyIeNqP6XEznJzAsSIaRsQd+8EDOmSOtAdQNQI8cOHNjbXisv4JD7lCBtA8E4g
GszjJBY50ziP8QVyf4/TtzgegQgZRehbfjB0HHl/uAoiCf2S6kiELxPqV0fS1DaHP5fTz7ApvufM
S7iYg6B0rdEvZptq/kMqm18uhfR5UUteD1AbRuKJjwPEZ3EokVbSulkbmpxFOj3L8XwrY1t7lIGz
S0Y3k7bL8cJ1j7bh/r1GHmEhaSFDgGIoaxWP2ke/DbKUqotglsB9iqcmnBTOi+1g2weQCyzaHLPi
0Aj4/qB0hrXVN/5fOm23Kozu6yKMNviZScPWJHOUlRdRyAoP7Tll84aW3JSQro2P1vXxFeYz2BMl
dt5aA/O2EfvjThfVPKOOpcRkPphWXAXH7GBn776xTWclChf7BuxYJP/F7JFUORHJAlBXaUJYJcgn
DsgMrM33JDlqudz9PtlzZpVuN+QoDzNFkY5AqbZry7bek2PJMClmjPWtFkvdkVyRwJBmaNJH/irz
NdWxhB9SZUJkGIK+GkCTZYGmzO5r5/JBTE+cId9khZ1852evJwk6m6tN+geprM2pNgFttLszenOR
emBK7uGsq5AtTs7dfsl7AsSUMJyaRBz1r46uq5yQZHbQN/Hi6OTUsRJzrQ+8rlapVh9SGtGg3Xrc
SkQd1nsGb5Kaha3OiL+kRPoXb//XzzEg7gLIg0bCsoKuQLNqGeiLVXbSl8d9X7LUOr0VcaBkq/I5
zE4HaXqzXDhtWNSvyQ/V7u7STM2vHs4lttaXmN4Vkr6qRSF6eoZyE11KVUbKuT0ApCKV06FStFyI
sJWKivLtKp6db57bXFwEyOlw2OKckY78hPySsqEQoRtK4bti+f5dLLfqIVX2XnFE+mq0p4J730Xi
KRDx7OhSdZlpAG4d1nbdLpIJ6zNgKc1ieFCoW3HNQxcVi0F8CUBGdB+DNlPeNa7dmcbTvM90u4tI
kAYucfeqLePoRobJ6t1R1C9KPpnG/bC3ajcnwRKyiScp3YEFiO8FfmKtEb+jDmwVYYY6216HHimZ
S6c3r8hBT1QLmcLyg/WDiPqI06qcTSGbr4yS0Do+tEbzg40Yxb5aEVDJHbAiv/bNW4hFSHgw6PP5
7wCqm0lrv+HDta+CMAIA3UdeLbvO2e5IuC8Yhe948s3BVaV77h/+fTtWIJaVN1akvbvFOnL1XnsZ
VW/dycOAn7ZGvOwTB3l6ilYcyu2h4zpITUVQdNrX7HVWVqPZUXb6+PwUjXoUqXAq/jbzfq87Wlwg
5d9ojIKnn8Aa2m1z79jh6dSvD4Z17S+wp5AEmM+FH2AsGZotSkf81s0VefUZvM6H+CNjnbvJ+KEE
07ZX3j9dZOinZGWCoUuHZ8tjlftC7mxc0jBKWnmcTMfJTD1mVoEBWLJlzTCHdeVgHpVr89YAbUrj
F5iZo93IAiOqovyezlM0zPil+kA7nMPgnXUZi0g5vV5aNJ8Cwgu7EQzKq20gw8JaLD5JWT44APQH
IY2SfL/5wWtGQ/msCO3H8QkpLTE63VHtXOUM4N0eIRneyMHfZuGbor29VRpyH0MxwHPReMUcgXWL
UyDpPR1rel76oVwjTCvLrN1zSxhlAPCXvZfqL8FK+YSepaPjSc8sWdQRk/+/fdujQkaFfPWSAaZO
GbDRmwNp3U34ziSGMdFbPpXgZQl6S34+vldw2vsQj1tJkaUJiPctzJdrcVPErtuox6joCS+siQK5
i789Xfml/zCAsHaj1v5FA5thudPDJfRFEL2wQPnawgH0zniJnurOMI/l9vDZYGIQezYcfaKdcmXy
R2b2kzAJ55P7alJbDLQjuIewOD3lwJUFJzs5Hltv7zsvjuWC0j+5Fg2PlwB2Y0JOx3LqTQE5FU3D
huZqb/s5wRvYMstMdSzt2zSjZvxJK5yb7ZwjbFEoQ/oTtCGsi/N57P0bAMizDLdltz4gdWiBLyS1
Xi9LKKq1vi13uRLyWyQcqFRRkXp1J/8JY8GhySQe/JtT4KchfyUjUbLskup1F8kfUddXFALdfslj
g31oHjagKRiWR2SFfns7ZJXgj0X+YkwDyjGxj2r/r+GxpCDd0LAqY1hLD52ZUlkjwsFC6pAOEtx6
vR2qu6hKpAJ8+qKlk8ylwYiAUniQdsQ3B3MwO/lRcK2DBFqZg+T9xSF1ZRFQv7ygDW3Zu8SWrlf/
Q9Hou+EXJ1yz+egvD33VurBuYgAqG/ti9n0tvohWqcUus0OVfZZ+u28xd8XcfGz5Rwl2jdj6L/FM
tfePPXr6Rz6PyNTte1L2G69gJ3P8FsBLx/qJnSjCvrke8CHbp+lRJUkAn/PfMjtpZGX/07PITU6d
qvN/ihMcXHBeH1k4AHV/bQpmom16etnDtIwagvWeEM+GNs1P/tkkbiLhsvMNLJFVbSJ0yj8sUoI8
VHTkfbIBPvDcENrCyyQ88hnNJJ3KG/UEHMgkUnCzQDWa7cjyAShqv4XEw7MrKpaw3aZk3Q4KfP3m
3lBj8eUxbwg3PQYV1WNH2kQ9OC0A0AkVVTsUcFkNR29NmG/ZDvxI1RFf0W9KAi5S99s+rM7fzHAU
6nXi+iKwre0NU/gnR7OsZO89CwNcArw5E1UaYK4mEIBNbpvUZd8Eq1/ZNKPEYZST6RJgmhJ4g5Fv
74VipGwFmCzibCA9a8kACHDsUNaGfN0VZ5lrfiyac0hIm0r5UrvtRdGjZkNtZ5aO4rYSGM80RqUN
y1hRagqE7MUMzfahKul6/oDkcYOuLpiUcLkgeYXzdgSP51vln+4K8gdEButKmO5I+Ua4Fi+QTYGT
n+x0kd1bu7MChG9BXD6OqeDi+ul3KOs7WPD6OShgn0BZTA7JWxlwjLXfys2Yz5HJNzmky5JpJwam
hFBwsd0D+DW/89ag8H8LiP96Z3McqWyQPJI9kWRlAoK8Al4YsRN15iYYACKdbwWvCITI7VONCS6C
olE8K4QKCd9enD02P6ElVUI47L3/bcQTpVYpiUxjvPHDbp7DBB+Cwx9XQIK7uFgwPyivt7dx/XvM
v68emUAf0DyKh2Y7AF5Tde9JgyXLlERP/6LCMvvXFiOfUmMfcZGvhjZ3xtkdeTJUHLp8ZVSKAKl1
R7cMxV+AJ5UbxZAp50HpgmdOTmXcDUsQ+MQqR4H1as8hFBorUJMm
`protect end_protected
