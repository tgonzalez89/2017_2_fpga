-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
1bUvotQRvcltxZDxqAi2QhNKDN97QgIyHBOcWH8567/wCe8hM+ymuwFfBktDy+h6RFMGgMWTIxpB
FpymLqm1s46Yf85888E11WeByESzbjc30xKZImiEp3tSlSpHYzRN/7BjcPA094X6R4PmrrPd45uK
VomRAr9dCujnxJaHPnXT7SBGRNzVnDx4kSyT8jv78miJmH2mJmEZ1mQGPKMoprUMk0Xi97yV7PTb
yhW1Xb0HDuCVVScGNInfCDkU4mpGm33XMR5IIh9lmF18M9eRDTYGXZMpdOyJrZp0/7/4RsTeitm8
oPMy2i6ngIFKnZ0KPh1A9yMEDP+lH/tHgSxuRw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4544)
`protect data_block
QgaFL4u/nvSdFRjcA3Uwxd1iFzL/YMYthgqiJAxwGW0FJDHxagbU0cMU/D/WwKSgzg+0fiVo7/XJ
nA3cv1Dr0VMwWATmwjL1Bqqn+TAHpatNMRjTBesaKfulcgA2nqbOrjfBhYjo5qmghRwFAAmsbkKQ
159gd+VovMSgKUvVUZM6l+w3/KrKTuA/qqjMWUm8v0sbfQSs3btOTt6pIVgeuTtrPSVzcicrLIXz
6cGGfVrHHy+rKMA7SF3yyNI2Q+Gk9lxufCdUClDkuTGbBSLjURB18d1wZu6IWMEHPbnUYp/+T7TM
vS5Xeakyr2FMFQ5cEkF34rppnt051CrA/Lf/qg0DltcznGu20gnNSbkjzskI5qm9vL+7bIW/y8Eq
WeBf62HMOHXzv1MUPhBTa3a4rn0XsNXrIOYCTUojjjNm+k2kvET1jrezpSNu/epD+kJO1yRjhN+m
7XRISVJrT8URYZ/VT9SKTw9Sehsirak0RAsn6/OV/6hTxKAefy4rbGnFMJlCFZVyHFLcgCss2Mfz
fDW3+7lFjOXcN6GdF867YhzMMP4ZcdtgvV0RpBmoTKNXqWQBo6d2jBb6C/m312ygutloEchGTBnG
APiSdfoll4AxYk7+6LVvagNWTHQCoYC/RB6XdoUurRKwZ4vgkyYg8ZusBBr+POX2CqtMMi8uKOAl
i7PWkjMMudaRQEYt2CXS3DvlF5IzjAXr9ITrZfEybmpqVHzBcvdOUBm8hJ89SmrkkYxo827foz1q
qNkcl+xk5Gu4lHllDW+QuaklkYaXJzEE3GpDxyMKPjriEAenSk4JMXYCATfO4g0PqyBLR2DuB+q1
C3cpLFIc5x5AJ26uIj3uJmBVFFJxCZBEHlPr4jAiPBMvXmtWzBpuhE5/YNkm5Gp8TW+rP7kgzyF1
aVcwgakMltJp4qiFHiJBvt2qfaUPB+DFktcsXAMJaEP8oYWRU4X7i5BUI9Uz5f2CW2kB1nqUcd/Q
QxlKErHpGpVjNHmaplUvHldGIZEjVzOm1FafRPUXVnKwr0dVPKZ5LA0sGBENWiwxmx4pFPbYEopK
hdVefUSdD+0NDLzcQPcLTr0Yqluw13RzGnagbEAzVKjJtHlU7SSI6H11TBaaIGvheg9M/n8BgtjE
yywU3JWMeDy0amfifuvoVMOdtdOGZ7qtdZrx08283xfx4j3s8vGRAJ66V+ka1bDjib7nENYjgjUI
ipp8nE7EfUHVbggpQxjDVXTvXNkk7G0gA/RFykRASkr4KbXHuTfGTu7N6OB3JUWA7NEI/ML9ajpE
0UMHCq66Hh1QoiCOvL+ME+m+cIz0WRIg9NRigIrwAgSwCV9DC+ofsRIcVXsxnBCsrwawRfGBJHgX
S0QyLWftb9JiG7g/U3RYOJqkiV6etZWCoFWyGL0Mcmn/RhS8GPsxFM7HfgX5fxuTUmL61yRC8jZy
SobrbYoKhER2RhebjN0CZp9b9dbvzaq46lcHCp/oBGmvId/Rv9W6RhkQEKWj/EkvFopmHv1tOyvJ
z9+GYCKOyujask/RLJwOKP7/7cPvoXnHq4NWhbnnNr8S85GbUJ6ySWvqugVxtr6scanHiWezBImY
b8atSyUm2yiNbmjJplofUuhEaDW+4CLG91/TYIWTwL30sbYT4+1BM68psEKEs4JBcmW4HvMEHOoD
fpicrfb2c6xfauxbLxjXoWW1fTZqX8KyjDR3L/zxZoGSEltYMtZ63lo4ZNvxLnrB9IyDEEKaJvDT
FkL0AsHstgwnX/Sx/Kcubc5hs1SAZMbF5lAScS8KXzIiKkxxVKmbAWEv9U/MPgzg8qZivAK0UWHy
lkLqC9mAnldFZwyi89QSaLOnsYuO8NxpRUcyrQgMhct99vSESF4hympYBVZ3mjg4h6Q9BUzgzvrE
HC4oX+PrbhDuw1EE8LxCq2yiPQSa2jeQvVCHjLAuuRrqrkqjuMCpfTtHnpHYHZ3V4W2eIyCGqkel
wKaJ0+/CGLcjC02HJclElpoY8q1yDDY0iTgSeRSM2XmSE1hRrphChaqHQZ+iq+Kfvg6qUbmerGxs
HB/l6HS9sD1n4M09QpZj/JM+seTazhEfxavaV0E6lR521bMLJiuMf9BVOs7YtDTGe/txKDiCb0h4
MQjfPfJO8HtHzKbzMkc83R8IMqMJMusdPxerBThsVwXjgyWDEbwERQER088LXcDTxdAVf06XGGwY
LQt5nIjfEI4fYMiQWV+wXfg7QFVFNsCOQrKFwOZHQmeoHiR63A+AW8HVBqBzUn1y3kfKBkRihqPh
Dwy9zdTAy36LY3itConMAfEDR+jgWRHY8pcX184JiofXxmLc+cRC1YCCYIHBYLKVIc856Bd4/UzD
PJdJ2rp6y9S8OB0yXGjQWpGF5q1Vg/lMuE5IiXL0PAE/7gMrRfYccFlVlBDpo74yeSKtOlWbp4b0
Uv0UnRv/7Zf1HUjMkdOkJ2lrOmvX4NAi6+T0pnQoyzdUExClbfMyFo0wciqdJFz5L2kIqOuivvN0
Iro2+fBnxTpmNjuRIZ/ywyL5CYwFMFqrQ39JvuhOnbZC/dHHRr5eRiQ5+0s+eDcpz3aGdByKWXnm
5jn8LIejBA0Ros05XVc1plg0hZlLiAe3C5L7sdT63YWh9ZEgPnnsGEyn0f3AyIJ9vitVUYzi2u68
mmhtqT1D8m2IBtKnEPpstmvRR6cIAWWHSNuXrTp9dsIsucgyItzHKS9fDgHe9FtquCebj0lKPj6C
LnzKUr1jm3rMeSMFgUChilGuGjd4dGwveajogyFeqfnF4xY5ctsO1zp9REaoxTX9f7vTVnpJjPYd
S8905/QJ997K4HIIzvjDYjjmSuaoA+OjMVF9cNomFUonKqu6JGazlGqLNsSwrmTvc80kE4HQXZ+a
bGUFpLao8IC51RA++tksfJATF/8n4L+1iRgvI1V8Xh0MX+Vxy2v2iGCy7N3c92ry6/LgMtypdHYy
PPrCG8dHkDwevqfMGjNWLCT+HniwJPHB24uNTVM8T/+oVDH3Fv6lwdgJrIFJwy4lAfB7H2JydxNj
CwkrP+/bPj5qkLLsUsY0u8TDZoPuyG169HdCEAZ3l1Vbfmdp9OVnC455R3u+TKcU4YJlD1XzLgfG
b52PJzveKwfHM58RkTFTI776xoeUVn2PEk4YSyJJ546JyoHHyB6Afo1Hj+HH84GXzb9ouIbCK6Tp
9q5UMP6wRTDmSk/a9h9k88Ozn49PXVV7DEipme+tB5REXRIz5VObhoXpWSSwCz3UZ677rcGR3BI8
kLbO0BLH53E1PtaKogTqbn/rev2xbW5yzdBqKD5KnfejT0Rc+1bsxey4o4zGiNWvaO+zm/7BQXQD
G9pUMg91SbjsEeCABS5y6Af8BbPtQiqZ+AmabV2IdYzu7dZHQqqgxI/iQNCYigc0wh3xkk0NUGb8
3Q2xT+uhOwmVlWB+eBSqzku9QsVs+QyAnK49kPWCnTBuQQ9iNQMXdjA3o8ca6eu9d36qWYdQ2jRz
yyPv0jTv3LRq995w9Rl2uRNwIXQQjbnYG8TXZAG8G1bln/UXjrxRHTup7QCBOxrK8PuZGT2tlpJm
IvWn523Tndv5CdcTXRov9Mc+XZOsVBjRkN3bMab/mBwh9gEmmtDUYFhsz1s/LEt8Yzi7BSQceYK/
pdwxlvYmQ/4XnITM63kdGd8NuxRwj5CJ7mffZKoD64cvDG5dTHu6zzoZcTFmfmAI8ijose+EnsT4
KjpCr+5EVTmPXxAbqYkoVwdveyAbXjF24XAm76FQZz7492XZAoWijvGMOlJ73bRttdxv8Xxy2Yuu
3+q33CqS/05EzGwRkuFhN3vAkblJfm9Lf+VEXJEWRK3rGnV41/cHO1bJnqRicY+eVHuksvbxdd9x
qdwU8ZQ0iGnRMtwBf5sHoQ3GZ1z2Kvp60bS9fFZlr/gNMXSzd7xuavS5RNN9C3s6UZWdmq8beOkd
rBuJOQGCKyOseBFV3bUL+sGMqnczkRq0VKjfYMO1ORQr4ni6U4xKlsDMgLo/Dk/FZ+K+hOCuZdEq
JZwVQtS2jvv/SyNyQE92+VlmSpFz139N1/pB0M5FIFDII5rTim+sq3xjYvCbP+7Y+5fWndyg9MYW
0o65NwaiREy58y6pPyXmqBmCfJrQjX3sR6+/QlH0E/TgzCNk1kljp4ArTImvJuqOVK4g2QRUxa3X
Kpkhgq9hYa2VMf//T8K20dEICBb3lGmwSPCsuIk4MvMYxQdPm7FdClFFPkyA8tQBUbYAGhA3BAb+
DDq88VNJO0AxRQqQWpeVJJcRKl92hNxZ+/w9JaYxzOOPFWI4g97GZV09JDpx4tgCZ+ZgFWBm0EdL
a1csJQLAl/p/QPp/yWW4vY3dBnSadupJJi13hHaCW4FQNku0HscUaadpmcsiBqqSbwv2aWujjiTE
oaOhPYpfJJzY4F8YfRc7mcQ4AwWlxVlMdA7gTJ2ssRyLvTjSGLupaujlwJq2f5MqzV5QgfWuMPE8
L/eqchRptvscb3Gm+vZDpLkBQncnR+UpB1pY3dIpYCuToZfTzp3qvLdptu+fRNVCOZyIG4VNIPIq
9ZyEP1FZmEM0WtzG84SceprTVrKIjyO9TIY4DnJMLIzsNkdCY/yHHCQKQSnlDvwjjeyPz+m6U2mO
fs+8mtRDfe1YBd3ReZlZt5O5HPg8ZwrmAfJ6qSYxzFkqPLWe/9JnuAhLkLHVSsLgJ2bqYp1+DEvW
XeHuNG8t2f0B5Wdp1LlXP/YZmiqpiZ71vG6YYEOmOZIz/0xuCdubc9ae90zE2wjAFE1QNMJ3bgw1
LS0D37zd3ut01NomtaYuWg2jxS3eH9V4PuGTuGScUFyNpuMY6ZGst5S6U6YhMOPdnh8RNDjFXvYr
4fIiAYoVXm/QIwk0Fg+TznoSN75T0zdOs0iKNAZT+hiN4QttqDjfTpw+AmPnksPU/F+ao9z+/yRr
Zn2hHgPRHddykeApwUL1ecuggtSDJPDv1TzYk7ysiqcGAWszA9+SJi0DSsMc352DMsHW1IfganAI
F8NpDxPGDehj77g9av+gCZkuJJzbubZlBJl5LPUYm9d+wEmKX0GaeTYuWrO0ZFn9u7MVg9DsekiX
cQz+3TM+E2Gsm+6pP+WHdozZy/sUHnrjBAc8a7rFVP/NM5TuSm1+/T5j4IXN1UXZe58qAHpRvu50
ZfugDTnT0XgUHzNQWWRP2XIIUh8SQnKjgs2/bd/28kosOtMp8oElV3bYIHi4fDNP1glppZidV3uJ
8BIsnvwGRGDoqehjB+qMfPI60TM3WljJVp5EwDEaW6sdfKygs20L56JEEDhPG+Ffj/DCgXPgb8cq
35JBerO6Lk7K3tRjcs1twGlcl9y+HMYHtmX8YJ2q5zYcISZWRlNTqskDZJBVTZLw1xpW4KWfiP5V
5/KSofJQ/jx/cIpnXnJzzbqk2jHFx/I7QufsWn8QpfOP5v4qyNL9qqWhX2y0lWokJCFAM5xUdSiJ
tLqnLUMVFbRAF8N5t2L0JFvqRu567CftA4yvVkYjhwBYRPMw6p+BINYHcFo3Nx9Azx1hDvd8LgNM
1FAuqBTTNZPEOeLOZoHStOILE/iRzYNmlTWfOtaVV4TYhK8SMEVvf+Hk4piXAWauQjHCAI018t70
xLpulsemJEE4PNb0ivZwDUf8Sgqa1oMAl6FpU12s301QbxLbX5Gljg0pMxNNT+3V3jHlmgQeCX5r
eNdJU+rcpedPy4INpylRqhRaGWNmw5IMsHLKyiHFpwklc9gqiOeXHl6Pctcv83+MGP3r35gteOsg
t0+lx8zvGrzpy1eHb/nje3UHDLBqyXaoLcRbflHodc1vQc1wicX6nbXu45VxUZ2H8cdNZMFnQVmp
69OVGVtEG6sGNnpjQWXOCt4WhSctf7bke4X6rv1T9ibpmdcK4QtLqkcksWhC66qM3TdsgIMpocEK
8tk8HzFXxH8iqZtq45GudMKKhJXebbpUrdh1bhDKnXkTcTBFuJiJTXtNYVOjS2yZdA3AeJ5xvWCc
S6jTQ/BZ87+KsJp9Ou4aT8XqePea59xd+ef8l7oiRGeMwVylSQV2lFU=
`protect end_protected
