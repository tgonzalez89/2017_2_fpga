��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR���[{�T���CK��TC,���:�
&��d!��]9�'D`�"9 S%�aQ�`!�6������V�W�l�a锦E(�\gC�slu�4U5=1�N�m��l�9ў��P���B�@+yg��=�}|֦���ָJ���P�P];4#g��������ZQ�*�J�T2�V�X���[��W�C��.��F�)\���ELԈ˕ݛG��\m�`iH�|r�˚��b��[֗ߔ\�z�	�e���Y��|\\̥Z7�1�uY}J���l��݌�ϑ�~I�3g�����E���M��������Ȭ-�
��k�ܬ�;���B��j�Ð�h���2�����uw�MXȇv����l�] ��._(T�nL�v��O�5�n�;�7D��T,u^d�Ҏ��0�v����g�uT������<oc�[���Iyưu��#�s!�]�e������),�S7��F�/zݸ���w׿Y>�L�(��K���|g+*n���]gv�H<'x
#��v��w�$��$i!�\�l����V݇�^zAkQT;~����f����>L� ����m��tN��#��o��#�D#�	N��H�H*�8VYƑ��ؔ2��˿Qp����� ��v;����98a��0�`#���j�X*�{�����IE�ԫ�%�.Aɣ>K@��rm8��9��K/* #���}�-��H��u���&yrܲ�S����3��-J�6��TΚ��^C����\�F�2���m�'�P[B;60\kK��%$�b�Obq*.�}��X�2�H+�y���]�Q�S�^���B�;���--76�<cT<jr��]��RC�PB��"N���𳝴�`z%�X�beuV���\�<�x�Z��D���|/����Q�������kew�c[���&ۍ<�1�*s�~j�4�jL+}#ЪX�rv��r�LЙ�Ot���BH�՞l��?�?x��ϗ��}��o
<$g��A�Z��,��&���@6j�,d@�8���@$M��"}���Al!W"���O�kh��n8C/	�Bu�"�Tн�YKb6b�g3t�k(��tL5�j���e�L�B+�9ǀ����ƽ��(C�=�=���� ���LW��o��$�$���"|s2c��@�@h�/�N�Y�z0iV�&<�X��j%�A�e�=�Գ��*Z
��&	������ �.Y�������������}�&�{�H�Z�T/�� _�~���Ё}���x���*M�m�)_��!2%Y�(A��zE�lEG�v}R)]&d���!tg�K0��/^[?���#I_Бp�|J�B��K�rOn!����k+z�/��V��&Ş�Nz�s���#�	ֳ��$P�6���+��lR�/C�ԡ��=��U�Ht�(`���b��숢(���A�h�*�͛tv������~�@3ۈRm�a�(u3-�NhP?U#�X;�X���RI��0�	n:�bsC���vs�X���0�%�N��>n]F�9�WV@1�R��3�ʇ�;����VX�)�����#���T��:F�Ͱ��原�B)bHG�+'�� d=<�=��g�T�y�o/훃t��GP/����_3�^�E��n&�7����Gw��&�5�_G��P�Y�_�
q��%�/��dTA1Ɠ��p����б�Z���9:�o������$�g�xۏ��?�Ө$%a%��%/�F�O�� U�kA�G�/*���Dh��6*�r@5��r�c�kչ�( �U�u��>���9t��-8ⶠ�zIj�N�KR�Sc,I�X'�"!�5�����R��"�g���Q+�3���tҚ6؎neX����E|��O{��%��)�wy� S��i5�|�I���!ʉ��SNR;���%�>��z����U�ˈ�Vt�g ��+|J��I,�i1Ms�����G�5�S5te�4��M�#���� %\:�K�(���ȗt���ʄW����l"�t�R�����W��zR�%2i��Feb�^�������Ԍ"���$����@eחքN��8C�X�F�3L��>���|S���H��e���=�u����8FD� �dH�{�9�ԎM�cpt�h���% >YrqPџ��Ӣ}��k&|�M|>A֣�f*����{ӽFy��4E�ٍ9m,MR�E>�	�?����FB�^����侀�q���x���z��/�7II��!:�2�fi>�He�ۏCe�0Z�J��,�<"��R��ȤC\�pY�?�$ϲ���� �;���Ͻ�Wa!۳V���j�P�^��&P��H�_?��臇QX�f �Me�x`Q�H�c��s�R��;�5����(���Ͷ~����7C��
 8;J�#+]�*2�~�W;b��x�:&X��T�N~yof`�Cz���ڵ	N!�9�/��i����^)l�1H.�����3&Q3�S�:v�s�����#V4Nk��${�m�_w�л���O_^�ni$q��h�/]V�����c�}��!Q9�߈}n���.;�������]?���1�DߔnK��,KG_���6��n$Po��]<f�����
�q�����A�28���[��d,}6��_<���w7Ǥ�آBB�R�O.�"�R�K�����ck߯�D��2����������t�	��:HV֥9�H�_}�cʯk��]��̵�a�hH��TQ�H?�h��D�[���h� ����Z�=��}g�n�����~N׃{�.�? �/
i��w��|�Z��`�;�G�a.A1g%bS �u�A�@�����*�XLF<�"�x��R�(�e:Z�`���X�E�̛�+A�K��,�24�Z3Wo֪]���:"r�k�grb��j���~�	{TÄ��|�.��2>�Õ�1\O��t�d��G�����)|�m+�u �)V @�*��t#XQB.e���!y�r����jÒ�z�H��xߛ?� �ge��pRq!��MZ�I߸y�cЏ�%�$��=�˅�����8`��	>})����C9�m�f����pH���@=�8����)��̺:`d
 �ǘQ���yN�	c�A6� �MY����7<�"�%�6�Ϸ�;��Te����E��V&�_����S�RC����D��T�@ü�fw��8�T�NM���f(�#*���>\��/�� K��1�\SKQ$'��;k����e�.�4�o�����߃�諚[u\����G�=���ծ �����Hd�ֽ���Y[̌��\��R��p��4��m����d�g�M
�1�B��S�h����/A�R�,M��t�%"T��t�z��9>m�=Mg��S܎�}��+7�߃��s\n���zoG���s�Vv�W��Vn�=�\{C�0��#L^3\E�F��ZK[c���$�^�k��]�vQ��ư�ↇ�_�E��o�m��od�A���H�$�Sΰ	�m�^��q�L�{�E�?>�[� �
9Oy��=�K��6`�<|M]h�����U:Ƽ�粋�He��J�8�2�#����a�]#��?���ަ!!�:���/ݩy�y�i���l*��-so��>�1𳮅Z��*'�#�II1y��N��=Nz�2�(|;g%�{�sH o�>�e[mh�P1luh*w��4%K�`e�@[no��@��9����\%�CH�AMmZ�����-���A�|��<0�&���jI7�����]rH-�UM�K���n�
<�}��/�*,�HZG5~ V�w�CG| ��;�2��T�����C�ݺ8p�;�x��7J�+uݥ���BM	s� w�&��!L���tl9��M�V�-�Z�8<0�D7�U\ �Y�I��Q�GT�@r�����}.���g��V0�ֱ���56����·c~��[�,l�;�*��j�'����K�ý�8uU�$6<��KY�HM�OFk�7�K��b*�i_&e~��ȏ�xt�Vw^U�x�,��	�Q���{s������f}��~�,����ҍiX%I����q�V����3�K�x$v��p|���Y8\��c��U77u��þ&xD#����;LR����2����cΧ�Pu�P4�c.��ZW�\Mu����N��L~Z�L]�6.�1�VP��q{�?�C��9�0lhi���=x!�Q�'�F]:w
� �繿�XqO08	�{��r�t���ae�Qu�d�";�Y�gK}��­W����H����A3G ��g��!h��?��dH�Y|�2h�8*�~�4o�}d�t�'Xw�; w�y���� 	x�&~�h�-�ߛ��Z��=�w�eaXQx}��2V�/�,^��N�	��ܐ��TS6��R-N�[A~�]�H���E�d�%���W����~]��/�s�k��� �_��5o��ؘh����u6)R혲�c�o/�x��6{����[���ۯ泗/�ۮ� ��)� ]�jnOһ�$��Q*�����g�H�c�3�}1���J�6&�ș$6@cT/�ʮ�����K+O#/h��pk`JD�e�w)1%JME<ل#Z*�lI}�kp�<���2	~z2��/]��n��;�X��(����D�%OIz6O��^��>7��E,��f�5��4w���(�jd�&j��Bu��#�z9���D�l�6i��Tb֩	�+F�b{��վspDe(���CK���|�ꑘ��mA�f�Op��a��'�����0�����k%f��D�K��x��Ēh����Izx�3��r�n6-ħ�jO(�y�{���:p4�����q��Ж���Qy������S�\"j����=�͏i�>�2qņ�Ǣ͛�^ls_����9vǙ�Ă�2����9ؠ�y(4H��&9����F���9b`,��0ٯPz�`�X��-d���/�0W��o�|JX��	���Jo1|'����T���D�}��̜&#�H`���H��8�;��Ɛʊ"�����rH{�ί�穙���7��c�eމ�C��Sa������zOZM�nG�US?�*�����l`9ۙ�3��%Mso[����^q��2��D����땴hy���{Xc6�S|�;V����v������1���7���U6-m�>y1 ���@��;��L����d1P���i�%��lY�����x�|�|�F�NUL��<lf�P�!.C�m7
,8���~}����z�v�z`�meږ4�o�D�ߛ�]��$�6��k�L�<��iT�;|��f�G�����O�`U߾��f�{��J|��iT-	��4m�UwZ��T,L ^xX[[���I���-���1����vkU�N-&dX;Gr'�Lg�B�G��o'F��Bxw���.EX)�(�����F�Yq�O��N´,4�P�@3��R~V`��}�&ึN��\�`IZ��aR�!<H�>>��M��\t[$}�T��Ɯs՚$ 152vd���a
x�Bi���O7)4�Q�y��Ə����+.�� �B�@��o�uRڊ.�
�U�Y��HY��V*M�ï��p�?!�M=m��W����o4$w<V�?��@��iűgy�_0�Ԁ���zL�-�(��;�4P��i���?_�X�"t`�.*�L�{����WmX\10H���i�\����,���~<=W��Y ����oP�C���Z��L��M1��BM��{9�K�:����/b��tX}�i?U8��r-�^6@{�D��x&ܱ�hx2��Ӧ��� ����;�$��Z&�1�:9�����o �A\f� '��$��P�-�H�*V�|S3U�n$�v|�9�?,��-&�t�~4���|�[�V��]��ʉ:��Dg�Z�%U���%*6�]���_F�&�w�l|�d�ײ=��MQ��<�LuZ�@������(�s>⫿@�%l�JBiL�1Pd�jxQx��uk:��Lf4�)�'�~������['x����;n���[�O$Zu�:)�'���^s��'}ltFM��`�� �%�\z�ȹ�Z<�����%�G�����-A.*�K���s�8�\�'K�oК�6|��B<�Ox�]��cVT8�0�ŴAQ�*R�����~ý����g�z�Қ�(�j�j�#��Y8����"�*�}�n��`���gd���@�~���4�1�u0�຦�_T	��B���arι��e�������y��+Ӕ&_��k��B����>�j>ĩ� ���II�p�����k�n�	H7c�f�t�&�O��&Śփ �ͼ���o���UP�7xO=h�g�M��e����v����C���s�?�b��"9��z.�*%Ž
y�Ƣ	�L�5|�M'�F��*�(J���sp{�� 㡬�=@��T�j8Y �5�î�U(Y?VNR�#���Ϫ�4�ͭ�nG�B���V�������CO3ۍ����p[}2o@`�5m$Z��<���f�c�p��\�X`��a�WXX�H-���ْ�W�X������62u�T���
5���~���]�Z��#�o��X��׭i8��4�����cy@6�Y�ӝ���{���G3�|���x��c���k�W
 1<�֎�K�����r�����_q�k=b�T��]	���A
�sB+��>89I,}�G�I��;w0�m�YE��i�c�\���7��a�2�V�@�gø����,� ����:nηz��G�	h�7�<�z�_��:=��}.v���O���fʕ%��6�jn�����~�U��`�/���X�<���Zs�)��/G��OXM1p���N7@�b2�{�`h���֖7�&�~|�cdo�$���ڴhYl��<$��+Y��v��C�-�wT���y�R�s@�`����ξ�^�;ĭ*H�q/�#l���I�������LM~����=o��[iFb��w���[ʌJ����٦�J��c��s��L�1�w����R�b�r����!�����L���6G5�����6 <j��.i]�y$2�yD��i�s���������"n.�C$�v����2��e�����u�����N�����Ȃ-q)]�}�q�:̨%�<<{W߼l����.�i�̕�pɞ��T��<P��thc��vX��� >��z�Q,.3��:�Ǎ/	��V����X�k"��$$��F<@5L@olB��)o��%�@5�%q��J�$�25���-��D�+�3�9wo��a�|���ϐ�K��B�$<�ؓ�Ŀ<��/8�Hi��!W�_��)w�>7���S��7G�A��m��s;���8�x��n~�E�����HA���L���k�*� �N}|.�oנ�ef�`����Q���UK��Ё�~Y#�1��^
J��T�
�%�.�b.��4̙�瓠p�)�6_܎\�<��=֬P�ƖL{���*���T�3?�.��-*__`(�8\���XX!�~�.�����;<��}�:�V�F��r�Gz���gQڜBSՙ�Z�li���� *~<.���\�GJ��r$����
�,�ے�$��\Bt7���|�S{���6����3Rcb
jGEr`������e�ER�ܟ�����g:��!/��?X��PD��Ab���
}���: �M�5��[񶠅�7��jvs�cle͜����׬�("�4�f�x�X3_\�D3���*p�����u2z�ۃ2/�c�X �v*��{�!�=ݴx�t"��,0���SĻVxk-�N�>Z��]�2��d�t/�M�V_<(=�Tal�6K�58��n�A5#i
�I��y�?_���ޅ^*+�����g&���XEBW�rՂ��^�Rv0��9>���xTuD��"��q*����>�����e[�;S<�85�Y��BI'�9/�x3O�/2,�����O֜���;I
��������9/��I}�^�R�ua/on����$�x/�5W���L�IL�R���0�-���R'��ǋ����ΰ���n�ˑ�_q�!�)�R��	}���𠧨�J�<��t`?�Z�������|��D�ĒM�� A���s3�Ѿ2Yβ�Tږ���;� �$�����{DK�U�e��v]f�M�D��汕4�4��GW��_�E�����BY�V���RޫX�qヾ��{8���?G]�`��O��|!�4��i���*j����.7XKlf��`�\�m�A�X �� n��X�ΜHo\'.l� aK�s��>zȩ���6Y�I����u����rH��;-C0���u'�x섟ң�Xv�l��X3��`&�+j?��e\�Y"�^jx>��f�y�Lnx��dX�I��Dwb�/�0�0'Z�6��_�H�r���yT��mI�<��F:�Z���L/��?�A�JI�?I�k�YN�L���U� f�v%d���G�;Q@M^8�88t��Z(Y� �*s�@�4dB�.��l��cu��\'��2�#��ju4ځ�۶i!;����
�`��L��b�� j�9�� 3�BԬ�H*��i�`���"<;�q\��gV���s�OV��U��T9��4;ݨ0����q�)jXy��50 ���q���#��Ġ���Mt�܆�+��Ä� ��Oq����"BC2���9[�B^k�+qs���1�~q��}"����Q��}�WqV����,��ݏ��X���5��H���ܪ�����;�#� LM #_��o���w�t�7a�E��0jϘ���!��jjl���G��Lǌ,�}���`L���δ�A�)�å���J��s�Dk��"�Bj��Le�|<���Q�-&�o�:
�v����ӭlI�u!b^�zX10�U�'���U�H6�_ ���q����"��u�����TR��V�/R�;Ƣ�yT�/�^����a���y&Ѥ�~P��x����&�y�9p��!�T2;��gQ	��N���e�CL�"��8f3���ߨ	���y�25�M*�~g�y�X�L�.!��0*�AHؗ��!0��@o!6���D~�����e/�B������}!����x�����9рAZ�&�����}��w�T�2Mi���[8���9��8$��p�D+��z�?̷d��I��0z$�6�;���<��@�m��P�<I�y���0�)֯�v/фr�[���D�Wj[�ejn��7�>+�aL����J��<1��C}E�Zd��&� !���i���R��)�t���&��[~�����T�
SY����-!�k����q-|��
\��y�|����P��Z�p����A�/U{��-ND5�H"؄�+����Qp���B����U���1����\ټa�mj>v�0ę�����۫5Ou��9���3���<i`0�<\�O�s��ޕ�{�	w��y�7`�P:8�B�8�C� �V#ڷ���	�;��t��y8ڳ�)�aL�
���g�2�t�����?�>�/2���Ef�B�Է>��3�@}M�;L!#4|�5���Gʇy˞��Lb6�������/�R�X��l?��
aB�����ې{���]��Vw��N�Y%�l�dAp4I�lU��x䦬<lU��L���D�+g����3]@���73�; �\FN��dc�O��v���"3�{��N�Pq=9�"��~F$奎-��ȋ`�
�q�e���H���X�m?p(�'D���3L�Ć��u+�=�_�0�$�髧�}�^y��z�c�\�@V�xl�|��qͤ!T,���@#��#����$�����V�9�����>�ܵ��Fmn��q��(8#����d�s��LN���%4O�M��#��4������ql�������kPH��G�j	u5d$g�4-����%��N.-�<�Z�����;#ÜP���������(q��ld��ʐ��1��?��V���t�dljUQ�qk�Mvw1�5���i�=�'�I`��`S�5U*|Z3�C�*}Z�&����ӕ����1�Y���7-"o[d�*j�a��"0�i��B
Ɣ���5.�h�
��ʯ���K�y? d5J�7X4�Ry;��BWd5ˢ,o|���Ԟ����PX?kX��Ѝ5ڵњlܦ��4S]z�;�M���Y�~�]F�yd�n���m�I}D����D��V�f�:2@�@cq�lϽs�K�NX���^s���K����x�N�fbÁ������h,^�x"쓘������X��j� 2?ok�Ҋ6���Ux�^�፞���{�"�*e0`BG���u�[��ƥ��ȿ0d��,�2���#��x0�x&����L�)�m�����?+��L��	W��y>��l7�=g���>ݴ�N<���F�:t��������C`�f(R���^4�֘u�U9�'�~�8<ϱ��{�&�ˊmjFl����,@O�R z���pG3<�F�))c�����I�c Ba�t�K�4��)�̈́Tb��F���߀�wH�|�Ug^����RB0��}��ƙ{2`eB��C:86�����i��BD�>$�5��ڍ���|�1q�6��@�m��;���'���:���nP�i�_Td���'��z�d?������Q^B�Q^(�Ȟ�F�K��c|��7^tY�7�M��er��;��]X�Z���?�=���8��6��H�s�qC��,)�� V|Cl�{�l��
Tm�͍��	�Iӕe��u祇v8�2�t�6��I?����ED�ҵ��c�P����4[F��G��#��D��F=<)���ث��'�C��?R�옘b�����1s�D�p����$���w�$ �]�Hn���7�"x���ؐ6�2B���S	���Ĵw��~u�t<A��*�&��Iet3D�2 8�~�+�h*�;a�E��P1���V7Ðv����|�����̫!�ޒ�N�����4ş�q�6��l��D�:ZڥB;����e9E��k3�g��*?ͳ��eE�yw��.�1S���8a�AUp�|�pt��b�)[��Yy�l����Z"j\�W&�dl��
�Z+��1����0�"��ved��.��pF
ȉ&��<�7s���eۄ���|���ѤLF9��k�<�d���1m�0�qabc�i�)b�`�r�AR���M�A+�I�zQ��^�w\�/G0�+�ڲ���s��`���ݢa��b���]��En��f�W�'h�+��gr��0S�"r)q�����^�K��Vxoۃ>���C��֎���R��A���v�3��n�x�-a��N/;�p�{"��~�#B2�p�8@�:�:�|)���d�ԉ�n���:N�����Œ�4��6��PQu�耉]:[�n)I?c&;u��|^�����^45iĿک���)'Fxa�DB�/ʦnt"��3��-A���LwI��"+g!PE����e6�ޤ��J/��7(j��m���:�q�/	V� ���J-r�%23J�4�!wӜ�PW�b.1U��n	'��h��*h���}cA�ǟ����0po�V+y�>:8'�O0�h��i�yZr]ҿ�y��?���i��_=��K3�LX��c40B��������2�>�fL9K��|�����η��}���y��[���}�x�(3+������3E���n�5c{���W隗�W�a �I=:�e�kT���i�x��~o+BC� �3� ^Ń~�F�����p?����J^g�QM�>. d�շ��M�5��Z?2Ҙeњ�Ȑ:��>���O@.����U��	H��}�Bi@���19ac���+).�FM��]\���4㴘0�*�|���LJ����>Kb]H�F��i�Bͩ7}fx���/i��� ��'�{�S}��
&����(�g���y@��oGv>HMr�!��c"�)��eXX:ʬO��5n�$�����h��i��0�%6)#��{���<���<g��r��rPx�ҔX�bpC���EB��kŖ2��@^?۶�@��i��7�<&y�e�)�3�I,e� 5\׬2v�f��A@��뢞�Y�zi!��T�J'�iHD�ݚ.�������B���
��:'W�eݾ2�������15�:2ԁs������q��j �oI�S�dHG��eO��
�o�AZf3%*+��չr��D�	S��1���=A)^�n=ץ핲*DZ��Q�a���x�>��-*]6��P�� � �6i�ϫ�+��Ƶ��D^��X[�7��UPέx/m9OYJ�y͜\~x	����v��N����$��1��D ��A��g�  X��P�(��b�z��]{�u�̝k��k�N5
������Q�ݼ��=�䞈�fo��F�`��Y�s�o@M�v\�"�5���qx���+�Wx;@�Ͷ���-;!��$���=>��f#�4�e�D��V��]?s�E2��7Va�kͦ�~�L�i��i�%dpi�
}'��q�w���.6bĲ�='���n¡ �v��n�G1��I;,M��l�nNd9�$GE}4�L���_�Wo�i��Z��߃�6��4<�$/��]�WR��|Q�xJ���j1B����05	��ߕ��q�.(o4JU���*h}��Q�Ch����Y����OޗTSS����U�*]9�
�	d*/�F�1�����;�SE�&�
s]���a��|� �e!�����j(��&�t��(����ԋ�-/խ���H�1c�L�����;��#�rV\���O/�3(`��\�e��`�g_��L�<����lة�K��s�<�LDc1e�"��� 9��mqj����`�����N��c��p�T;� �w����Dz���bD�U�D�Β����f��+��͂���{���Vu�;��j67���{Q��A��P���E�T`�b�)�����lu�T� K������|f[y��6�+����6\ ��e<�ěq��y��a��'+�<#Wà�������h�C�
�E}�h�p��Ɣ�DT����+}���{�J@z�����mԊU�<v\!g�Akd��D+aE�W��V��s+O���������y����v+�I�l�����qe%�B�ŗe��8v���lW������G �`A����f�AJ!#X��L��,/f�T&�d�o�?͆0�f����KP��A[�Xe���ya�N��rʎw��ڔ�ɶ!^�h�&|>w�~�мت|c�΍�Z�	Z����̤r��U��� ��
v=���l"T-�y{9�
;�!Ӹ�n�i/m������ɹ����~���Y�NRvO�R�}�-� �����^nV����~�|��~px���ũ�&sa�Q����0\�<L���*�� �.���$Qo	�6Yñ�;]!��L��2��<�}�u�'hG�n�wk/��_Y���V�'��u��9�I�>	�F-0G�fz�v��7v)c��b�;�"���=��A��>��T�4��b?���Y�{V��V����胤����[~^Kyr񄲹�d#{H�6StV��+�߷����<��s56��?�0��oV��,�R�'N�(,{{�������]U^����(r��]�˱':��<GjzUc�/�u�����s��r�T��aB��?�//Kn�Z�_�������"������4��̾q�-D)�v9\�js�wg�Ȟ�+����X� S<�$ot��r#/lJ�?�m��)ċ��C��,耹QO�-���y�g�*��W)�M߷y��{~��_�CbB�TD��~�	ch-���/"�����j<')���Tj���?�Ut ��-��
����I3ݲ~[�8_]�L%�����7lLŴ����WK��-#읢���Р��lȶ`6|�]$�6�����9o�YSQ�&|�O���
_�ZI��US
:����?�CCO�Z1������ &-����JY(.q44:��
jyiAn� v wmo}�Fe@�#Ybc �����V��~^!�ϞbNc�{�ꡁ�3=�ѕ�V�H_d�nÝt�b�HG:h����4Z  �aiͣ��̽�8k�����J�;Ƴ��#�գ;�jd0V}
9�)h�Ͽ������+<t���SlgU�����Ikv
862����6���;�������5�ȘI�;����JD�	�H!�����в�]�LU�ܔ��%h�A"|g�_[^l�����8ZJ	�k�AC����R���D�	�G6�KF����"�g�M����|l����/����hC@׶.;���i��sڕ����E��NE�	���m7�Z��B�Aj�**X�{{c$iyy�6�4{o*Ίw~���F������*�qFJ���}[�9��Y�V��!�LX���X�y*� �F��'�RI�T��a���_*�P�{pry_k���z卽����!���Ԍ��m�Z��>VyB�wf!�y���:��:��ӿ�	�J���i�C���E%�&�m�p�q�e�T(R���
."�e��S�������RmR���ەB���@w�p���� \A�i��Կ�د�U����V�sS�/�
`��|���#�xd� �5���-�Dy��7�:ZAҮ0|�,��d�b��``�\>%ON�0��������FM��4��r��H ���ђ 9��KP���yQ]�S�ǡ��x��ݦ�V�8<	��>�qd(s}�g��aT���}��ϝT+]�2#̅���Uv�5��m>~��썖+y �'amaS�vYs�.s��� $��l76��H��yz���JE�4Bw�*�N"�t@*���ͽ|[0����H�ŗ�!=g�X�h,�ݨ�g"8!P�V�E��m����n$���8���r�뛀�#���9��l?��	&��_,�-�jΎ��X�����\
E�*�w0����a��N_c��f+����*�����>Ej�Aσ*t\A�&{¬l���۲��1��E�i\/�1��0=���U����^=�7��\i� T��n�$M���I��g�	������ ���@-���H���q�#���DD�M�Z��;+��a��ޕ}�G��F8(/�؂(�Q�-�f��p��U_[y?�;����0���J\� .��L+"�j�k��p[�;h�ծk�7	�ђ�� c���QC�C$~b���2؞�A�c�3� �J:eB\E��|/�� m���%�v=ᢀt�_��WZ�^�P���+0�c1��^J��(2l�B����j�f��S�
�.��aUE��t&Fc�.zО�
�c�4�=Ss.DJ��1ϛ$��������t����ґ鼝�T�R�2�y���9jX�~N���C!��ޏ1m�!Iq0H��/��":}�j��Gb��D�[@_؈,c�X��1�A�*���(�����ޭ��\���"3>Y������H�cTgg`Y�s��ީxм�D����E؅#Ϸ5�_�c5$^s��@����|��wS��q�����(.<��zx`�G�;�=Ab�f�x�"�L��4Q�K9p����^d�<H^�j֤��l6r�T�F���A��\�! �x��lrE�,7�D���:�3�n_�W�z����P���N0������`�x���5��f3�����6_y�y&qyZr[�d����J�.�jz轆�����l��%!�p�\���7���m��>I>"�@�e�����;P����ՈQ�:��^�핯�K8a����ڙ���;Z�s���)����1pU�������K�L�	�?vn�j��M#s��r�@bP�d�SI?��
��,�nGsײ`���صN��
�F�K��Md�w��p�b'�f�frN���I���GAr��Fץ��Ւ��������+�5h�1ŢX�_�ȋ&�I��feܒ�3A�X��d7��1�l�c�B���å2x��2gE#��IF�T��/��r�m�\��̓ z�٢J�{��D&��ښq�.$𞌍B�-PD��dA�|��2��*(	Y��m3m��xs��.�0�x�H�YU����㱫LT��%��/[O XA���re��?�����7�\��1���,C�Ft�h�^[��\y��bp���-G߼$���������!)vG�ŶYtd�.���6�_T8����M��bL��t2߶$1��8 ������\M4��I�6<��#�	i����2Q���_G�L�4�,#F�j�rK͹1��gϵ��7V�ZI�n�Y)��T��D̓M��gF��m�wԫoD�)o�׽x����\���~�BVm��#�L>+���kA=��^��樂q=2J;]�m�Az/�s�O{*S��<@U'ې%"#�{Ȅ���C���ϼ~��oE��z>˾)��b](O����xg�N�L�N󏉫��c�9�|S�[�S�*�)#�H&���3q�͗ e��U�L���'��YlG�`�I�_)p�z��@�T��޷8aO~<k\��h
T��fG �/Œh �:���#��)f�x���>$�,�A��g/��I�uk~dX���J
�щY��֋ueq k�,��+������X;`E�M,��ˤ��e���)����B.i^���G1��ͬ��\~�(Ҝ�NjӘ1و�HeI� �ywr��)�B�s� ��}�6�Ca$ �=d��c	��2b^���&��β|��4CG����>���7Ȓ�Q�X��B^���� �Z�E0 m`;��5K�Ra���t�f]E��+�/OH��ϱ0�0����������,�Ag|���ƚF���������6�K?�W �К�B�W2�$ԁ�!J�.hʄ��I�}�%ޛ�w\��#����Q}shv�k��.di��g��zjHR���
��K#���'ᘰAx W�.�/�����#���K/�f�#�9`[gי{Q�49�J�c�~���a�������|Hpz�V�g!���
�bJ���_���nj�J�%y�U$�t�YI��J)X�]�$ё��{�g�~�IM\A? '�(k���6��J&4a�c�w3���KK��IJ�h�?v�`/�p�망�������W~"R��eq��2$���.�窓��;KŶ�μ-��L��Յ�C��2g�dlĥkb@�t_Q>[���'{��T����am��x�*�Rf]�śT�e�-B�l|S{���Q�G���yV��g�pp|�=�AAU]�6�y޻��Ў4�*�V�������*��j�|���"���cx�� �nA����W���x~e�l`�!�����w�N���g�x 8?��J"v���X�m7baI&�%��B�>�y5��$�6':�UN5���<4t�}��@��P�o�7��������B�-��j�yt��AЎM�6���Wʜ�(MS���ZT�D]h�bF��R��B�Z��	k*��V�0��̡����2���ʼT� �^f�	�YYd�S	����\Ur�.�ˑ1�/U�;;�W�8�{��eH꽕%$�G4?�St���Q&�@z�2���/�{��H�2Ǉϡ�m�`��I&����&��`	}v[֐���f+�U�xV�٘�y�Ħ�'_M�	��x�v��ChO�:+�֡�?��?�Y�>'����w����O�O�Č>�����L?xC/���{�b�"3hT��Ƙ���՛�=��?ɮ&n\S���t�.sZ�x2��i4]���i�D������������,�cQ�sZf&�񄗢��!7i>8���*��r�̟��zX>�,Qۗ�1@�z! ���+{��[F������B��Ǵ$���ڙXGz�4����C|{a� ��ݸ����SuO�N����,������4_�)���W�(����;T�X�!NL��u��]X�`:�H�k��Z9�[l�X���gRrBT�c��N�e�h���K�7���nMH'����l�q�%��5_�tU#`�ʍջ�'(Qw����pp�a���Bu�&cI^�G�},颯�jӐL[K~m4$E4�E�^I���bz��r�#����TٞR�E=��W�xq�m��K�<|{�^O���ޚ���F�z4�p��c�O�*�<�z[��fE�+[�����-4��U!X�l���_#��.P� k���#��ʠ(�Ks���wD����ڇ��4"ӆ��)��q���	���(�
mt��i�� �W���g9��A�r��Y���w"�v�S���؎Cv��[4*�[����F戧{�,�E��YB\E^��/���Qb�ٱ�u�c8�sx}z$#�{����p����ѦM�:\զ�P<N}���L�����a�Q�V�d�|��p��P`��j�^�$l�V@��+S��0T�覹����LǏ-Ο�;��H�NGn@=���3����������}<2C�kW��!+i�e���~뢾цSĒ�-�C
Ӥ�"V�Z:fж�)�r����<�:�	M�q;!��fO@�'2Ӌ�����]B�Oz �hjB5?�_��O�����:�_x�]m%;��5w�
��A�����Tj����M�2�g�Zqn��ʰh����.�}r[!��W��"kc�ғ������]>��N�l�����.\I��0�F�_ތҝ�e�H�l��+�l��(��H&.52ރ\�m�*�:�C��Z�Y�^P�_�.P'�B\"ta6�g����3r>nh�q�˶\���Y���=5ù���N�-��v�5���t���C�7����N�V)q2#�_zpcss���-:	{�}��d&�geפ��� Z�ՈH���yErfަߐ���_���"}��Z�!���dzM��L���Za�s�ҁ�C��b'� ��KX X�$�|�:|�rvN'�Ýxq���*.���rm���dC#�Q<-�p������j@��D��ӭ��6$AjV�ُ�8�>ɼ��T)G�� l΍٧~H����9�@��[�oDƟ����O1my���:��4��x'!xT��JQV�01a�&.����fx�s���}z�-�o�V��l���^)?��͆��i��G��>��HŁ�5��/P ��Q�����Xclv�_����9%3�)���t} �7� >pidp#�s{��,�g#k���CSQ�ّK�T&�3��v�
��8���Ui}$�(<p�Q}��#k�Iwk��cX'�J"�5�O�$�SO�p��zc	���D-\�Yq�&�s�z�Ҍ�}��MO�'�);sG#��\�vV��#=Tی��Xbq���]�@cG�|SB0�̎I�w�q������~�Dq�I4����j����?�/w	$����!�Xg�wĹ�y9M��s���e��c�����ǎ��]�E&g}.5O��)���(T0�4%��f���$�9��'�?ҵ��d��TnJB[�