// Proyecto4_qsys_tb.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module Proyecto4_qsys_tb (
	);

	wire    proyecto4_qsys_inst_clk_bfm_clk_clk;       // Proyecto4_qsys_inst_clk_bfm:clk -> [Proyecto4_qsys_inst:clk_clk, Proyecto4_qsys_inst_reset_bfm:clk]
	wire    proyecto4_qsys_inst_reset_bfm_reset_reset; // Proyecto4_qsys_inst_reset_bfm:reset -> Proyecto4_qsys_inst:reset_reset_n

	Proyecto4_qsys proyecto4_qsys_inst (
		.clk_clk       (proyecto4_qsys_inst_clk_bfm_clk_clk),       //   clk.clk
		.reset_reset_n (proyecto4_qsys_inst_reset_bfm_reset_reset)  // reset.reset_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) proyecto4_qsys_inst_clk_bfm (
		.clk (proyecto4_qsys_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) proyecto4_qsys_inst_reset_bfm (
		.reset (proyecto4_qsys_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (proyecto4_qsys_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
