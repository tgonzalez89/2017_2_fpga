-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Z7QpxGGDU34Cs6uo167yKu3NBkDJTMhBlx6aI3eEB3iNPINnHXo8vPi8lXT9glsFQw9QlXtQVwgj
/B3/lKq7zvkMAL78mTpzhwfhGuSiDta8dLGlBTwjalzxbeX2oX7/BU41PE95eGKZurasPcLVj8JE
W0A9WnRnIoDn35tIwJvHPrcU0lHgllQsBQIfXsfi100DO9aLORToSqUraOhZIFbroiCqoi7yMukc
Fue1fuv21XbePSwynh1v2IBW+CUYQ828V1vxyC41mzI37cznOCsaeu4YmTXCN9cEs/vbIR9u5WFD
1LkSqyJvAkYhxLBuc+3PWRcVUG23DPR4X+qwxg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 114048)
`protect data_block
p4eBzztMXrZICXUGy7qRLurFhWyCab1u+LsW7qp2AaV3AHLPH+4gYpZVypwSSMB4LWlHop1DYxFr
QCTST9UFvYdOVmlYlJab7wsGz9TiLwweWCKLKUonpywLhGtusUMylifWCHOcpQHBuRK1zHXXXLYw
1h+vwmim7uMCS7R7cPEOcZNlnblvHp1pwJ/3dyruvVWzdQfKfowpGtHWJDmd9rovBpkeXGvmSiqU
VO9m99OTcAdR0U3TlkoDtxXrPYOkgeLtKRGhK14QuPyMGJVehJIF7q/pXrt09cyJjpV+2OfUEQBi
7EQTh5uAz6qXLffeP11bsedx2t/hInMdZoPMPeQC6gjfuYv+6uGVP51p7PhU8VG3T7LeBT/VryXs
elCsU9Oq9Pe/qZjlAs18MP4e9WyZLai1Xssw2omZ6zjy+g/6Xg+q1DKu7Yp1RwniNC0GV8/iMcVR
pooQpGdyvtNN3HNch/uE+BRMfRLFu3woMag6c4+Uq52PzXzjDzF7dJ8FGEF2zXWCjsUvhS9koi3f
qGGbGqxn1O1w89V2Hz452P+r3F8wV2Ojix//QZwWefa/ZE45NNdEqmVl/yB6jIvRpvqYnGf6fYK3
MfJIqqSCSjXEHIEkrDag/s8tXYjJdsGKC2X5qMKvh+wtyLNRCN2fmtf4FYII27a6Y2BjH8yT0nHH
6VRAxNrb/suBnhRT9yfjQmHFePEEigJAEfv4Uw4xVFcmKdQFQt0W4+9ab2hP7gKHqqW1XjvqjeNO
Nf1EKCKb+zaCt8fHsLiEysCW4YSrpT9Ph5RLBd/W3LI0H8DN8ncnzEm/CPrmjjP0VxTy35yhImo4
+s7XT45HrnakZKiFqMSmUW5L/1yJJgwyChcJ+PKyTbl812K041gh2iG1/CHca5u4HR/1XDD+oJTM
FILzJ4upV3OQF4LS3b6k6wZPn4WtJNkCuX9shmsEZPgUiQgQut8TO9A0qoQ+sLSjhcySUTGJqIuQ
7uYoX25tlcw+t5LSzoWXf0O4zq3e5G1UcMzoiiVwiwqtwCaiTahJLfGG7HII3dA9wOWuhNZYh4PZ
7BrYVjYaqkoBu1Rb5wL/zq3+emhc4aJ3q2t+2HBwsBcSqBD+XEOgS219HeaFcEgDlxDcIPZh+FhS
ohb4qJju70/Bm2mYZI60/nwQIa2DlPJG3sFRFeQK6UkKiiUvWgH7h+cGJoPfkSIkthmiNVcy39it
XMUq/en86iZKzlukUaNOh0hPhXdmqjfyqn3IXIPfcnw372zedYnOcJUaMEePkA83xyHBBPHhmAoT
OlpbJfqtdVQ+mfZNxCA6L1R/kNsVYJys9mGiReF0p9jbHWO2Zi1iyIPpLFOfGDYr4nq3V44hGHkO
GNvROOgtDDF2e9o1WUgMFpFaNVnr9MW3Nfd9yg4r/WjqPKMUtbQJv+KeFxnWaqeFMnxiguOKICrl
GBeOZj0Rb+2Ga0yoV3x+EWwm/cmFk5A44ujpQOEsx1lPtaqg65BvBOy33j+qHy00noH1EDaPqz2E
nJ12MR0gfI5n5lVZXI0ruHw+f4u340ooqce4D1SSSD2MFpJ7quT8ZKrGaVjZDQFayWoN5w/33QaF
Ceo/m/HEAB7q8PgMtpJJb+0Kjcdej4QTCF2pzqN7zWSQMx/NBMv9hrg4nYO6NNy4Un3tFzCApbcK
ptB42g22BT3Q/fTZwa04y1yyGdts/Byhk6ckA1/zUv35jJl//j3RhI8ipLDeFQ0vsKJZS9TXY3tA
nE3Uii7qTGKCHR10OoxjVRHwn5Hm1v9Op9WYZ+fyvdf2WXbDvOfIBgPx7BOWV5l/UcuJsqKwml4z
q7tBPmGlWedzuKoRniFZ81zqVVJgZ812tizH09omTOEy8Fc6+tXNcZAFYGfd7FKb2a03GYzkMz6H
iQLy0jEt6U8rS8R9+9OORvF6M7cOmxqL+iIIDiAxmnKax3IQ1ETS/hStONZdqTi5IPkTSVFWIQcB
rKfPvrqXAUmF+EZqVXYwZi9HYuyLljOlY4QcHUO1MmWzS/xFBC8OgMKGV/xSsynxLEmvyxsTycRx
RL7ax7tWqE7rMENEn9eL+zXkE4Ogghu+pNjRoLDRuLMzaXNNDczmXQ25xs5W5gW54rc5OupqpVEM
LK6EaLo8pY6AD4Nv+pDXa0gvvoX2OkEsEIK8AKoblbak18GmfmNrI+Uk1aoHOZHYkwsg/zZQLOBN
TwEQEr5Pbd/dCmU9vXqtut/DWAkgv8BeXq+s0C0N1/UMxZc6gDXvsLjNdHCChQzO5+GaCjqtnoU7
w0sjFsLVGQ03htccL3cY2ZhgZk3cjB2yPuFTnxBrBeP65uSN9Ov1nqMYtcE3XbV4Kd4ROPstqhY5
kTQtBYem+nQc6BSrweDDIHutyHcw5Zm9JbDx6NL46GoJg7Ca4CJMmdn3MpXmhgBl9UBJCNDLNK1s
EOwNdxVrxx+Oj0YGssA6e9m67cIeo85CmPfQBh+9T3e4JKgA0iF7Obh9z27t5CODuRGFXqtty0vI
MFoYr5pwMn4Tb1Hj3GB6ZSBNmab/Vizo4sbJtTHoZb2t0VxLXjOEO2yfWaseYAFSoPr0F9QWKxLp
QCJpQDr5BBXyilaEGuIHCqBdrR3Dt1r+Gf+2QkcIgWUFcoFqyMn1cs0qGktCtsKIY5U+YceGCGmY
3zaXqHOjxneLqzs0yYEmUx3famV7BEclU/Sj3skUe+fHMTU/DLYCx3B9eweMndX+iCezQhxFVC/o
6HNOo9mJ20n1d9jxVbWGnoVeP37Ue18hyFgGdlBHf1Z58INDhAAqmRY0Bgy+7Ik1q+U0PmbEz42P
QLNqG8htxMTsY0OO8VzBwouql1pjEyXfIC4ryeGy55CxrdjbZIce+NZ5AzcHtQbPTMkAOIxL80ed
FyaV2JcimeFGq/IH9Z8+6ZlARziLxj26YL1UdSb9CQtW9QBFjqCkIz4QR2REcwfqNs7tZR3jjotw
LS9rC7iduf3mHkAs6mbTIwBkWkTZV4jdqszwO8hcB3bliAP8z5B+HWCVI+Ft7f5FPHjhcgezr/GU
qLzSDiTN9h8LsXFQBgMMb3zvtmiBwpk3BbS8fFty+gAtyScNdUSR+ZgcXfVQt1E6Q73kbrUUZloc
G5se/BnEx79pqnt4xWuD+JTEX1Oo7JVc6NkewD4fbLZ+g7sIsaE/VcEfg9Qc9MHbTYU1+Sq+ThyX
NKElbJY6D8A+/tJ2NncC3lJ6FKNWHTuSSfPrlQP0+Tl+DAwWXOy67CjQj0NSBHTPnmIjLIKP/cEb
vwyletusr8/EVhPpcvid1JVutT4B25AYX7oRems5eY2Q2g7m53suRv+xY+D+pYiSzVxlT6cDLG2Z
VQQ0h2YTeYfacCJQFjxVp83G512AXrM4qu3jEsDoqa05nPfb/31hwKlvCy50RxR5V1n2iDxdvQXk
QUmIzd36XN3E+BKsMvMHb+zf8UpE6cypNo+WOZM0Faj89BtwkpHbGjDJ9EPCB1Oai2PJemJ8Oxy4
taEIwcEIssPr1QSlDM00MuGFIoZF0IxwYfT6g45vYJYsJdGpi5pqFOa7fs3iHTxRDIH3d44yPIi2
ZCVSte5t5i5ZM/GPv2oKF2GYFd2Y4Dpqf6Ljj2bVc2zgk0qV9roMfMBsPu0XlWTaEXEsv5TQLWa0
tZImyI3UheyppIY/EkfUKWrYMye7qPqBBO5pzhMIg3hy9qebpvBwikcC51dbHi2e/z48aMTA5ACS
OaQ6NEsYFLWxKGV+Pm8ibRflcDf+hM/9iONN082Zy3EMD02mdw0FhXXsoESS7sEz5nI7TdGH6P4i
AypqC78MaKqU0JcZVPVmufwf+c4JBek5zfN3W2eNZ9mC3wNnwkb6FcCGgKIUOlE3Spj7hz64gH4y
QUQCuH7uHy0wgARQMsJoffA1ky/4VPmC1Msb4iIUclWRWOoz7LP5gLreTpa3697PnZs6xJ06fT2w
2JSgE+l0OiRpP49NjxNpXTqtm1agOdDMW4Gn0l7SI6vqp9JDcWGxGWHkioufWbavsEEDsyAj1/pc
AEV2p3fGHxG11jTFduaCKJ2kcKhAuw7gr1T+lqHFsFm1uu3gDHIXWW/stEnF+EitLUI8sb1vLVt1
ARDmfTLMOnkdesHM0Tp5x/g8rOCEsTz5oD3gGGhKe4eGeHabwI9xTmxFl/wv4xh8ca0zuYOHoGlp
koReS+xcgJUQ1ZU8i+vRAogp4aa+TlK5OjwqR4vh/xTc+5fK1MUIa4TSAZ5+2C93EPXqIuCn5lC0
bRCpEmzPxdt3GA3QEUkPr/Hs4/mcyenkSeZa/PS6Lj8j4hu++V8NOyuwjj3XFQVK2BjRQGCj8j6f
jxMmewsz0J+2q6CwWG0/0ckhzlAQ7ktmJUKqbLl5w2L/Tiy6Y/bSCod9NnThRlV+HsfjTQ9ziS2/
NHiTt0myGj1mItZFLHlwZrE/6kvuboNW4cp3nj5oJDYDTwCvVnlwHYhtbBNYPh7szPpRiwfusjRk
q/TSSowllrLOvFguDsMzV+uZn3arGlQXF0eN2L0Y83fgLUXpSX/D1WKvxwqRqb1sJkP6AzdP7eQO
ChO95YIeAT7uj6DL/Fv02WNdqMmaGmk1agUHLRgtmEVenpZp1/NHJq3VIXUBLg3FslgicNTB+sVN
OUxGuVJrv4SyxCMXQ+2ktXYrKqqUuJAypUNVZlqUxh9mXr9akivb/3z5/vsyRjQqYq18NPeziBu8
7uk3YHhcUTbFGmY4JG7EDqglqWXHvc+ROdLsrziMTfoKBMFUY9pE/Mw/0VglOs+Z/i633SM01IJs
Kw2RiFq51U0a4zTOEJZc5nt8TPorysnAu8f2FVHEJH75sFcO137I7veHblCHr8HeWg/DT+M5YQCe
ucLiOsN6XqEr7LnJ8F9vqH5PW/p8otvpA+Ed2vqmteVuf6NkhAAUwBKA9TMRqmvEuRn0oy8I4Esw
24C8IYsXi+Ow/h1Xzocyjrioa6olRvQ4Hvxe1uMx4HBiwZu0vdny/z1/NIo1brKGgOgd0VKq2NM0
IhInBk+BjsQOK8/6BM5xWfsFs3iig3LUSneprSZJbmeBJdqcJyeD40zh1HaHQCbeGmvboXfdO2Hw
xd/PRJ+rco09MGhSSCclD/alVDFMUY7289pzXAuKxUYBJVxKzCM1w/cy/TOtv36QitUtGa1jAQjZ
/s5hfHkDgkcTmndLyL4UngxAbV75erDAPi9pDRMHD0KmnLJlR8zHiY4dyN3Q+IIBhkKJ4kwcWYrn
lPmto5tf4unYP3s7djXSuR1NjN2z4hAgOknISfEFjJ2wVWWpF0Bs0NSE/qEFk8uuYYzz3JSGPlFf
kebk+OAQj1O94/NnoXhGBhqya1+gzgVlPZ+dUDrP4eW9eDvit7HzW+H56B+9kFYlB6XZqJCAIIBT
a8W2C2l9p+y/Mbt6zbf3tgDdkSJEPCqO0ORZREovbO/1kG114dvaKnunw4nhM4ei2LhDOLRu0Ybj
MukJK9TpnWi+rkt3uFPvr9iCHE4w1gMZaFtwSLyQYyWNSBUhfgZ6847Sfy8/xksohgBMmL8M1Gcp
Qdtn8rXsHpuUA9dGN328RdWWtorZQYPvsbFHuZX0Kw1CdrlqMqloSIH0JKtpgvSkg5HajCGHrQ+I
DlRVQK9fH2G79CuE0Qrt1aavQJmsdUf63Rc96BoqG/M4kHB5yY9PkuVuMjPFqEv2QUkW+LVJrl+2
JDH9E0vhwvjgJaKcjfafouQa1h1ZmrH+4obV8kKZw0xLEL5fbxaixDbgl6ZXpKF1uPFzrycsIEGj
Wqi+J6oAJ4fHZ01xfBnSH8VMZPSeE1Q586pUcpi434IEeDq7KkB8qefeDECOPt24nQP72RdQ/Jqu
ReMcNhIXX4GMh2rPlBv1kqUH8BsvVtDwL5pEd5qzHgimhVsB0zk56LkS6CBDJOFMPjz52q8Lt19w
NMdyJo8vw0/lqQLoNh+KOMxrdt+sr4w75T9zlJHFhruyB3SUNPdVTg+smoD/GGwMXrJKCSglEs6W
Ze5IAW8TCTO8WTZby5iRcbQxgD5Ivw0ZtxWInRt7wPXgLWBu/f1Xb2VDNuSV5HwydktYuabu83oD
qMj0KDqYFgd9qDJTiEGDkUImmv6klll7i9fmt6s0+sTUVuT5fUrkadiu3vlcXqMPmkL1zIYtE7am
3LKASIWyqbrm7rlrbQePNM+nRDsvoPWkouD3CnxLsGWNdzKa6YswwKK8ZKDcjS2ZD/CbMPu6MiLW
sDQJAtWUFK25Udb6+u/to6DTOw4yGP1NUmgjf81g3U73MbNiR/8ftk0MTkStupBEQ7HbX/cYyXuZ
eWOmAmkifw9DnrJexTXQfv9AS6ltt8yBZwZaRo4fCDli3GmhwTCzDZimJmErx4oYOgrmuR+NF0qR
hXmjw93cldqXt5RUBrSUEr7wg+mHWm8LMi0Gy+Frc1pQgCWBfPUzZ/3gbrgar7yn/yCedI97JbTi
udLTrJvTCmSFeFSOuZNEH8DDJ/ONe+cP5l9HWy2OUwoZfCKf380MsECC+FtE4cZv38npKGGec2C8
kf/ZYqi/PKVkLVk6WBd8v/7OOchIDT0rwGkIHa+qmRKe2aBrY9YGg36S/UIH7wxEHGx2IH2gfE9k
ewpOo1SMaljiX49dy7qMsFzGKk9AQ3hOU3OZsHdLLQgRLaFPkpgKy+HuJKD4rUy/L/x/9JTjUSXR
AjB/0eobmpCpNnPUOmQX7uQR8Z0TEsWRXFlr0p5Y1BkoPxwdiJN2Tqs7p5QP3zd7o/iA4MS+cPOL
+G+ga/mQ3G5leuSlRi0qvqK2k3dtAmC/UGSOPZTSpQ8I46dk4LKeqwjFMVaOg2aqLRdG0LzhJzB4
+bLdhaYGQd1cEw2l7rna1qlXA80ZJGOKjNrGpp0OsBeedgTNP0avwxt1EfBaH4nkZQ6iIhecsdO5
FCx9Ok2/f4ABfY5xPIwywlRf1OaX7hg8NkwjufY1L5tNALLsXsNdn3uwKubrzUTLpIupujqB/W3x
B4sTmt2l1bHFrvTw603kpTE4tWtsu2yEge6+sT8AFLq9g4AMv1e8/7695evW+8I++h7HQ02dKrn8
xxqh2W4HNsi29Pc+x+vhNPypH9BmEpbX7HyWsl78s/8yCi1At7FS9fOqmtroGOo6MRbYGe4wkgyq
2hoeMtaKcVoVpz00tWcjw+oUgkBjRPnC9a0uobRVN192mXY/JE+2ilXEhpan6jPkgMIzcW2uJm1V
t+TzWPDe29YnFaBuJQvzIMJNovJKU1YHnLpN+CfnC+9/9WqKXLoHVhE4ltomRGpGJnQqQJH7ySGV
X53CwEahWGY1CuEEFZWPe8RlYBb01ogFytC8FKGB6KbWZ89Mm7Dix9H/1BPUNJrP0ZR338XkAGdZ
H+QwzRxYXewakoGY8ucJVHR3CCeyyGxXE4QG/zyAQk6jOn2flEyN2FyX4/iiYmjTV0PPrMaEJSLg
x5cvRjaMJTRVQ6nIIGROUXlLs4C4Hl6ozrnrvizNF5zLY7RY99E7KGluc10NRwB/XuA7M1UmIhdn
/WARobeMUC6/ud+81yZr+CNi03QXfRuVqZ3LA7YX/bPI9X3/w3p6A5TPDc+zk8lJzpW0xuGCSGAZ
qRkboCpjwvWUXNJTKo08L7CuljxYYlpHpzKAhwPVdXsb1ogsSg1nHYK1YtUQYRJ25oW8Rct4nRGS
xO08J0anHbvs4zFcUNtUhcQIWBcJdc7CnAn8Sz04BHpWjPKWwzkGEvYbwZ2LHcPWsH/bKoKa8LB7
o+EUTaFXi9tl95G8LCbb+L+Dn8IQ/0vL3NTpCXblLNyzqQJTtqf9Yg/jGJmmiPTcinBeVwlsu+FE
j1NPvDEQOHGz66RFc+DvFhnvJIF9rP7t3y+ZE7/FojDQEwid3EjoxK4ZiGTd2aplFuyGFoUlZM0X
4dXaUjfHocA4q9mp/xSGSpk9BpMMrmJRQgZbaoTBwLvVKw9ZNjw7s04YQRQGd2lKRaUbauF0O9+p
uJikcbHHpl9yQ08dni36yQjqVc5eMgUvgzWhnQho0b0JHlfDHlOziHTg+Btdsi1MtLeDb4ovsV9u
CqsyS13BbYLIxdmXSQhW5vcMKPSethVfxZSe8oWYtIJFN5UUmETUveCYp0QDwrNWSEw827xXNB91
nDIK2alFpg8KQ6KH32rHfhbd0r1opZgrXmEKgOOtZkLJ5uyozCGOrUciDUKjx1dq2XrElY/qkhw2
O9Ehzm8DJCut/rHyimGPIBGLMHfL2BnEcVgb9toqzLjwjQ+azL5pYVShgPFtS2wD+zQfuXlmWxD1
MBXyqjbqNGGbyABPsu3MkmBVtPRm7Vt6JLtFrp6UvwoEyIVnAEGDuJEcOlixzZK5d5U8VS5fF3D7
rD5ndX4RLll0UoBipkNiwN42T/CIzPBa0OB2HtkUyEBm9Vc0RjZEVqYNusxeuwSqGnAucmzLSZ9y
kPEFJBentqEQxteJomd2OeedS/kVBgHt8lMnV1rES2t4opchF7TAXkzxdPXKAzdtR+rfpteindza
xcrMg8H+YVa0gzz26TdxFkXNvCaxHkLYs6+4BnSfURVGdkBzJihTm0dQUzBEoA/gg5AUyUGgClUx
i83RlxplJ6gxsx1O1q+ZBRWU6rvfaiJMw+fxyYBFGS3Y5b5XkxnFEq3HmKQMeDDTNdULgeHZHImS
Zbzd3KrmO6yQ5HfpO0a+rBj8dfvUjw/dzRXdpmfgY8rhuDsSDAZOtpq80plMMcAbYEVYJcYCPvQE
5i/u/9TG5AYZTPQ7orY/j0VM1Is/VDuB/vIvoIfLTck8jWZo1UFZieDgVhWvPikQzuzNJw5QKEpa
0foBUKuusPm3aqkD5byGp3NCyzcx2RMkEulvhCHXRJysQLKGCKTf68Ow5Sne5BQc/ZRzkJyBhupb
zf4L9v5h5UIMNorxoiMMl/8Q4jkD1KouRe3dJ1fWgT/mMzdTgMTFU9seYbo+uSef/MZ86wGSNJlH
JpjZWjGes5zvgIlopKb5GsgSpOGlmMYkatB3StxJ2VN0twhGRqY6NHrLdkmb6HBmZ1Q6/uYUAX3+
c54NqTwtrSaxFMcSuKk6CePK7iDZCjstNyjnoiswHadkKL2yjPEnjD9hL/semkKWe65kqphjdlpR
Y8AXZdaNk2akn3e4YUgP04JLBFnwX+1VUS4ZMRmENrYSbG7pKtutmLXHxsPrqWeVtm9g7Js7s9aj
IAge9/gzpjxM4kaYS3ShoVddPKkJhZLd9QCxt62QamS8W2igMJLx/kNm4+82SipRwMBpXz1BmErW
gb/2d+it3REGKz3UrVJItoT8JJ7rwXQ+hXfubP5rUEW8JLoyYRR7rXWMLOYBIMj6Kky9+5MelbcG
VFCL4EIxcD5br0WjNuoGmzVL3VP1kGqd4r6IoQ3gaZRL5ZM+XHOl4A5fKenBO5N6eADIiKCNkG51
R3Cc61k8WL+tx517lRb/xEY8mIKuWcX6nH5yPgPiICXUfIg6Ze6aRFkVtJq+/rzNkTA4F56Owj3a
XsXUdYF/KJ5iuP8fAXTVhNjyyF/ATgy/EjQgd2HA47/PPJk/874kKbwSpI58piKR7x2FzHpgwVYJ
fG79ul1W36RoPV/DDRBDDDeaIdy+xzcIwt+0h6nyS3nnnL5iX+G0plC3MA+ewYFA/4dnunnsH/mx
/DnS6/gztd8WdJZKvrPaGAFJUQe6I0FyaVdw2UsgwNb+WORT4NnjFW7JS64woK0ejS2YbKgdPWAj
Cp/hnLB3Uy0OxAuvFlWgDYfIpsQqz+dtOeXdo9tH5Fiu9wpdlOeJzjJLXeUyQm5/lFJg+TcJbMR4
4+hcbCtP89aOATUsg8dzHM1UaVQu1tC4DTRyJ3oA5KHF+xi/3xnfB2tNzJhRrSu+02vUkZvq5uUx
6xZRrmgec9OtMU2jIneAtkT3PY/32l9NFlzhSzRKyXpUc66XCQjWs+EuE/zhlAAUgeXDZHfxjy4U
qgYhgKCCRMCLjmvj3Tdz+k1hzKzdBZ3xTVLzSHLD/m4ofLEHmdYxz8T/xHNC/VWCEpv+0hOYL1IY
y7BVX2s6YJzRrlv+MxzT90rtVF9SduxtNG0yovMvbXnv/2DYQfpYBz7EZMDYN9C+nynuSFWT+wdV
YKbA4ocztvi1+5ImzUZ+7fvJShz7CT39msb5BHkNatagwT2zZtTS+y2L1UphqUVjb1e++MSrMMbY
zxZ355JeXrFOBc6anlZVwFTZZnSKqj7kPk2RbEZdrUYXLdSgDpivFeb5UoYFKls2x3byn4hCTERG
Hgu3fEvbIVYhxnZ5b7QtdpCszJ8KRcmB+kUkunR7XO38k/AarWG2H7GYS9kfCUKIPcuWBWm84jA7
aHUObRnufAJGL6eZ+aObEQtTD+1eQbOsoVw9BYqhMkBGdd+zxCvRCt7iWwyw6PW6STAZAt2W2ITH
/FqesPGIsW673Mxvdr4aGqaD/BRRQRUInGFEUFtDVsucGjfJDN0Ui8PQxwIcT9x/hGeFC5RdOlmo
PxexG0fXWxMD3oSHVfbON/HRVlXNsat8sHUmsg2YUFbamu6TX564H2rof5Wi0QYuipmxblcGusNa
F0yZA+Fca2nZD1j9yNykpTMbse9PVrVBu6t5nm2EEQ95yx+Y3eBiBBykfEh398+W9RPr320F9Rpq
tXg+Rq571/ACytcaet7qbfxcxkq1mCz3+6sWPMh25SENCdIzTGQjS21Yzw+qLawLCEJo7EzIMhUE
HY/v0esN4U1tLAmOAIByGeF+bJMEZVx6wxkJEWMP5S13FTO0m7RbD5WtvSjQInm0CWeD48HQUZRH
WT+o7frhnAePaA//1OnK02G6zsdSski3qj0vI3YetE680LYJiGuZ5JivpjjrzgCMaE5Kscdurf5v
SpX1+w9WxiLW3OLZP5lvQywNdtktMtzVbxD7tvaohlnrldFJsrcSJyqPjKMHB36fZBoH1gh9JHa3
pItE0nuhVdm9FwlvZDkEK5tS0xtW+xMT2N2vJuInexZUmnK5jLEdVQltoPM6R1JqaYshhValP+9P
f7Wn3ShpoFsuDQKaGMZHMqQ22WiC4Xui+fzaPyaOJ6QjG1/fj5MlBmnT8YBGw0qDTeBRnuVLZjmf
bklbJ4XkhmxbbiMVQ5yBKZr/qo0TbWqq+8mX2vY/Rr086OSqZ2H0JQ2LB74KFuaQuJdOX6bykf0z
L9z8Uwi5D2bnPHfKBAtQgZw2YPGhLGryGr8NW5wp3GYpszat7kIanlkVdMPA0n893DeojMC8T4H5
3HteVU0T3wf2FFSHhioYgWGwuL6BYvK5ZGgNEnYRq8jOhIcuQnQv/02jkVbndoHTAPJJu3ArYQut
16UEY2bkQ+nJdt51JEaqZZXUsiz3PAvEzrjkYkgyzhpzOUcFxb0HW6yDMY7Mz7RY2aN0yhs9dQhs
AtdW95UK0YP5hljdqStOyZe/qRn0S1fkr2VtD4Mkox67CMZjZ0jryfNffaI2omfdvBj4qJQ/pdFv
PkP0ibVQQa/1YNIzv0Oe1Dbuv8P7PzlAYZ8AuqPRs7HHWuseMZvlRS281lVl+SkB5RrAYKCpXQ5a
DcEPgIxyZ24CIuECyStPAS0Tf1GPbZ4zlzervVw2V3lA5UAniN9CWIPaJdJOsLiVKcwHYCVPvZXP
wRBriramgZraRXzMyd61t33I2Aa7TZ9dEzOzIA24S9tL2Jhg+5G+9uaIlcsme+NZ3JBCGniizi8L
y+lj7Eoxq5EQCNp1dIhB9qa/fWdaw3m+CZTv4osYO5SOy7QYsM/dTHAG/e08jNSLJgKCFZ/e6K+d
U5Cng/OqpjfoS7IPYtPPc2g+Rnx8jfLScWAHCLpAZS1SHh3DVqihJo0XLPpZzHVBCljXOadAoZ0Y
bJWWo9iSjz/E2HClyWbtv1thOyq/IQG3qAR74rfhE577dnrBncEBhFdrT1Bc9ucOTWoDlF8H0RxQ
76fU9bO8rz/4NH2ZtetGK1scJ17dqV6fIdpUCcQ1arrHvi7u4PpWqUMvvmj4gZp8EyOSUsItBEcD
r+MySqKXlUNQtK7d4KYcIkHo1DVz/2C7cNflSEXtrVQQGsWETY/bytbxBHZxlgVU3/3N5q8D1LxO
JrAruZistOVamE37aJKsW/YxJdd4p9LicAe5wNJ6RRzr0aCzYL7eRYBMhH/i9OuAyYJGP1OzsSeF
phsubxoGF4cxeFbnVGXDaTuXI6GwE7KFMUmAYMQDrhUQSwCEePswqKhT2OyiKhimmOU/lDouf/eD
/fysJmLRxATMtH58SxlibEHdEIf1jq3stSot8211J+R87a6mrO3PbiaIOh5qifdqUv570rLrfxVz
IQpisJ+XeJpXotraCI4wnUhC5BGn07IsEXwtZsyPgRih1U/iPuA9Qzfq+lR3bhFwv79IBjQTjlvm
/rCXmzbY1qaM8vbBjxwq2C0OogRUbwPqcBFTDNA6b0I50kVuMHNWIylHfoUHGK7C2eXBEeUscE2E
MV2l4wLvDokB1PnVhtCApTQ9ghvHK5GYTAYLn07H30alWZ323wAqa2XCNCY4eDkgvlkT05wUUFVn
SovXGSnxhhTJF5o+AxBj031t+8z0Ew/UKESQuzViZ4iqK47sYLpSsEITBzrJJ3FxDk5bjnQ767X0
14bcoCud+id6cs//cG3Yz9yd5PLq2snSiWByjeQUHljycd80f7j4DZkwgT2I4+y55o2S81Ej7vP6
dqwDyA/ksUzoGQXMjb+EAzM45uYI1GF/EX8/2iaiZsRXhtvGMzN+p5In7UVD48PNInT4jCHwxfM6
Wy1qf8l/SZ6fK84zmm74PKvoVaaH3nkd5ejoKlJICxxJz6MuPolU44YiHNIL7LuNS0cfqZSkyvaV
bLlxMs8kUewmnhq753/Op4gmpHYGYMzM8BfeYK6a138PR59kVDwmSYIUS7R3FIw9PZ/uQaaz9ZPB
S0uCYeuT8cSXdLX2FKoE6GBzk2ZvHKoMAZq+sQlcT8GmvM518zRVDKAl9GftZcQHXBVTCxOZNOY4
1pEv/pzFH96pPiKK6C4Gj8cggN0pH2FKQTdgHwaiqECC/RVx/LkPJ50tIkgG3YVs6i0C74ff2Xdm
oATJ1SaFs+r4lRVh6uXXJYb+fHIMwAmayABCs+WsBFk3X90hoy4Iu4Rv/czeJXhau7BHA31g8RVZ
RTNBirFSNudlbEj0aYfXOddF0BdaaG3jZTwIEtcHmrGqMk2ojtCJOTf/LpjLc51oYZZkg869TnLH
1gN6MRdOi8wigRrxK+2hH8Fz0kyYFE3YvlPmYlascErJp7sgW0w3i5bTrTeMKAIsCxFl/0kKZepy
f/RWTuxG0dgtH/050BC7XDVkweWucezh10kfDfw7zO4WabubIsnYMlzVxVU7zXNPA1Xhf5UOLG9X
Pulen3TQQC34ybx4vQIp91FdAWR2+FNqjKEdChLdmKY+9md2wMYXgkK0SoyF93yamTNTCliRbdt1
SsHyB31gNQeOeArlPolPU4zweTSXEDUepEbPclle7tua9yqtPfe9vSMCf1I42W+FLNXPjd0CH8WO
bRTSLWRuukj8sNoHiP8YmMp9bviT5NGGlvcyYME7jT2zk68SCHUz2eRvsWpu2++/hb4wvSXAxk0Y
OS/oFtJgKHJb1D8YaxPI69GTQltW2LcBd3doSOSGWbN7Pq+oSgZWwgH6iTLL+L56aAs0afskscQg
yYJ0lo6mTxgMt2EFKyNQjDFmm45cT7aGoFSvMp5edYu2CJ7hMO8/JXftR/9dzFboAkLXfIH/Ph+k
7UMeeVn1EekGFnHjP11eMaqkw2N9xeStx1TPK7dHOOUik+UCUVlD7ZkKPTEAkO5yJ/dWmYm4bKYv
YT/CZ6pLfMDvy9pwgmU4Bu4Nhbql6RZxS/Wwvz1lNiyIrj/OYFW0w357LxzU8cRojwfpqkjAnaSI
THQSjFgi9uV9TJqwh7km+V3JHsRnU5ljTwHFQ/onW2bzVJ4tznGdK5y/JJv2LmrVxDkRH5e/1/ni
8aO7lnA3Mi6XopY3MRppr3uIWc+KUTQ6hmE8ackkpIc78pOVnK6TUDzH4ItrPNIFRdyTSEQo/al+
LBBaACIEvZWXxIMFn9algzxZ3QmYZZGXnkBlD504oEOMUUytgW+PiReazIiuQqwVQQ59+qJI8I2f
TJo/ob4VOyhee/MHMoOCrtM5pbf8TqS7jA65GldTdCnxEllBoSY23HQQ3p4VAA4NfMEeFVAig5il
uFYbUBvoRw3gSlXb6pMjQspFEiLUmCpmMMMcinPUzjstm03mQIyxSbZnvI9eZuRsrsIBCE0iGAcZ
4NMWeC0EXcaLOFyjT4M392R9KljuZzBroDMkAju2p87yTkQKY6C7VqCaEHWjmNMykgzSm/iLPk7m
twDJBvbCJzVTHu7gOCQVkbvsBi0J1u6/TXV2nK3K3q2lFGGSbilDbsAnkvYAxR7PiCREI02TI8Td
ZaZW6i56J5ydtf1RsRtZThXRF/Mw5U3ZZy1UmdKxiKH66GC2E4bZq4tYqiEw0yRVPnLwDFHr+3sX
+ygU2BEHAncLoxRkbMit3sCTrYKRox/Gb7VUCuDRgyg98PGlJFhcmGXshLUooR5zrjBFm7wMHi4Y
FEl2TFaUZ/TjrAegJtuTWW3EHCkfHxDwx30y2m6NV0hHAkHd+A4wzPOcniP4x7NSNYFNIETRirOy
UxVU1f8l4Mds7WkeMBJdeQlbuiQMd5oJHt87n2+eL5iQCf8tigBeoXKJkE0swxJYLfilIvM7CvHH
7MGmlRyEMHIYRXsmYhTxpg5Dt+nCvaoSUWou0lYwYuKXhezu5oDzHJ/c2dOBLDYuPL8ieey/q2rj
wRUCJGMWAPUO8NU/60tdxADaDSSca+CQzngh2Fop/Qlzrzugwy1b1p4kcu6RGS2ifnRz3VXxYOlw
qbJkblDZSRyYoNd/8cacO0R89c1BK2tidSya+OzDCKcNws882Ro8kWX5IpYN4XMKcjK01+DHtJ4t
5hePErIJGvubRZ5dlieBXYiOBOOiVEX1/mbOI5FZKPHmzez1U6Zaw56+wsLTgiXYVH6wRchUe8lN
oWg2MoggfO5Q0hnYfeWs9CLLPKuAqSasS+7VcLOZ+qu61N9ZkCmewcN30kwpTAAIbjPYBPJsF7+W
ITjhb/RgkfXDVgDhf/6wPua3uBPOR6Fh5XYhdSM8BPbfvqsFTyj3G/dW7qF/tevYWsuxZU540Jpd
tMDwavyH5lmflRucYwzgFByGZV8mZG5urKJG/hC01unnK8MPkyTGppEjWykIH1dFNxNc8GGHrK6d
6R6O9fubTCRRiE3jU/lhFuPuKoL9eUBMn1B9TYY4Vlk8RGHVCty9062Pz2LmYcMyXrnRbhHXYyBX
JUbCFYd0I/mTi07ltmE8rpqQr2hCcKF0ROu9kxg//BoY88UtcXIkuwwP8UH4qXf03djRurtGBSfF
U1bCngo0kIMzQNEPI11K/9l7TtlMaqwMW3RK4lVKEljPgat8/vqnAv9nrMqGOWuRR1vBZSf+mE7+
cD1JnjBZK7L0znf3rWtiCnX26oJ9ixL9dJ0n+Nx8BLTDWVx2jsxYdyArcMrNlG4ja1PubEFKhBB/
DJSzRnH2pPdQCs8XeJgWKoEDTKzX+HNjzGi4FlnQyxAY+cMt3k9hC51UsWd6CxVWVRkixCulYesZ
rse0P1n2yqaLxbqBGENR733QIp1b+xjQKTiCAcJXatqd7g/V5bCv3CtxrqeYmDzBZf38kAD2X7WM
2Qb1GIlrbiUy+6pXg+fkOmvtM8Y/AVcyRDyQRcjC171bZfkHm0qULoRCYPLIWRe4G9J/iaP/s5jh
ybCSv4XaeN7atQh2sp8zNIATuEbnhMIrQCwup7qNoHkEsgaj5iSD4KUfXaf/woNRQGIv/y0tG56T
Iyra/vZeXsDsjIuafWP9FJhnYyDtTJB6fnUnKXu7a3W2c3rqv7VM9UGWKIZJq8+M3jJsaLqrM9NU
otsVjOWHYAjjsq13d1Z4JTyykwpKAZ1JfTOfUqWYLNpmEJynccQ2o+hFA7KqGkjj5be98fdew3Co
zJb/e5VkxXnPndUaYsuGP3PFI/TdZjnOtFSOO36BCHOUOoKRcLxI916Zobre9xChMTzlDCi6hlHY
s1Madmo8Rv6p8Gk6RjfCjlP/GfZN7dnHNnrZSZRNOzCW0V72TSoCByDMsHeFnOrPBPYpfrZwQdNq
eJk00metQ6aNpvYRK3Gl670eZkcPDk1xRtOGly1CVTRVgZCGiNxNNzMyPbcnUHeIrp7VYTiND7nt
a/W5COG+kxp8kysz7hpFneEqo1yW+8Bha6x1XTym8do7sbhgJ1cOaTKeBoMqBl+sfxMGefkCAv5d
oFGk5yosivbKTIYhzuk5Q8F9ADe/TWiuX9fU3babSPkctz6iQ8KKOR7R2VVDD8/BWst71DwtIKvT
HoGSngKiDujMn1rNLSBmve4NHSMqdAVpS24qQfUiXySYGQatG1TLg4beKKCEu4nm1kAmChYRg+z3
edxE2AJUDKj0BAaQTRN6bTl9v2bHm122IsjwxJKvjrSHNZJgYd+E34k152mHnIXhLbhSKcA+OM0T
PCjsNSXzM8KlJmbTYFSvQpntUjm986Vci3/nuOwYRfdKJ3Z/TEOI6mitgYvH/NLfNc7n/xp5fUC6
nPBRQTPCt/k5pNPIzn6V6LgeQsqBOM1fZMAb4qYNW303f4pY/RT//342I0ja7hmCgYbU89VZUEmt
SwyXn9Vc++lFyV9ZRe/7BntJ4jXeM62pYRoUA6Tob8XKAVrYuUKDpaQo3ZFfvhdsQetCDAswOzPM
2q5g0o/x7FFl7NLY+4KRM97UaRyDLw1ABH5m5jp7zFaMevDuvUX2rPzB/plqAvXnrg74Caf4E/ll
mNemwnruSKz7/WPqfvTr5ulnzm5IpFN8ycx8Gk41WVPRqRmk0cc4EV8P6vps9I3l2KGUeClgOk32
X80cJnIMYE1NCCH5GJbRu9wSy7LKDS+zsYAWQ3hxe/HIpHDqgnmCpF3wC04tHkVbeW5Wmfyeb6GA
GRCv5TsSNZpdimFZDnJhasVoOcXQgYXD71P1ULiINoU6Yr1tci/+wMDR7hLsP+EDXONIVOTzW7FN
KNBxO1ucr2emO73M9WmZKa17jUPRZSJgI1Z0wAWAMh3XS7lEhNqXAVV3xXbeN9r3c53A4zF0zxD1
+OHU4t+3ODmjKVel1i+HvKIA9ffZpBgCkZTzVHS7sFbsUrvr101/f9Re/4qFGdi83FS/Oczz/F7q
eu0hsla/FDocF7rq3+PtJMGAYRO/ddNelIgOOz4GEwaTrOc9/90LvFq4BdHSiJn1bxvihGL8gdNc
vtqxfxKlI4oYl+yPnSgs961023UEFz0lwlSA0krQvwSeBmkq8tfwbbD4Gjsqdva0TpRdJgpRawJk
beiDbon6Hk3pTytcRuabh7w7Qvh0tea7CuIkYzXYsEVai+yAoXjyd/PvZvpMN0Un1HWy2qYnOH5y
e78boujDTIuR7vx5IvgjnsgU9AD6yXAvuGz7gEmJt4gIMWZRbckqYKHuEEMB11Oj1xze6uBbBjjq
yDugIi7euqpL+zNZPKNjZa0S9cqtXL/cza6qDLHwQvLbs0f98JLS4qQRNSLfThkcLEfOTFwLsy40
LDZWwhDcp3JDS+K/I+8sRGZtPvoy1FSa7JBzG0jTkyEi9RIpo8H1a1TcYza53KgEAch6qDP5GMiJ
jW2Jc7FJEXisrAEZgbqQvzC35ROWg+k7WxQQa203UnIIrbHYefRSjiGtC5njIfCrw0FPouSiR4DH
B51DuWmpx1xmn7lvnkWhcJWqS6z+OKxabHF0nu69zFETdAd13JHsOsqIYLD4NAmPJJbQPQSoBvUL
Q+/eoHdbJi7fQt23cBcUNuSlnaHvDkkNc+edoeTNGApfZQWtljnN4ddyj+NTck+l51Lr78rFK9DE
Vmn4erk8Vbb+QH+BjN14I+SxG7Ttla79dRALQmU4W/alZwT8dJTz0OzNb3uCWd18YJUU21BR8HZI
JwNpKY20SrjCpdvSfxdexTY8byzPaMOco7gCNIPo+S+l6zshPFquIpeQLZZKh6CTJxZ6/+YL/Ppz
F9pDy/ehqyZ7p99ZEzeghH1cSfVhkhnD3SnwHKqZQRBeeuhesUVziLdCzE5kkcYYuzLeVWzGjazT
GkxcI4AMNHZ0S8Jm7JaakE9vEcwuVSmxnGJpYRq52QGypB8HIJ1JXZU/6es+cglTwycXzCTumQX9
oZZkqRGSfVaIeuNJZZtyt3v52VVi+zHGm2jpX1odKwV3f0ujgdBY8uo9IscytslqOJicjWqWiDi3
f7iUtzzQO3NYf0YoNL9H94CQtRgEcn1CoD1Xnlx+v8GBji6fQHR41ww37FELCh0joYPbBknqbDPU
2jkCs8EoMhZJIx9ul40oh7FVf7mhprghoFgwsu0LA5BYS6++N0annmBkOiwNGOc2H31Ejd58mbAE
Edxe3UfVLrrZWAdVdmXY/p4z7bBPdNMhTjvkMX5RcAeChmMZBom+ZV9jzeb5EhnGNJSa7nm4NpVy
v4VjmbgkHLmOwSQWfbyR8RRGbS83ciBLc3QE8rfJgULunPYdOB91a0Euh8fIYiIAdpjmifaAMo5g
vrUAp+quYfpL2RlFre2O1UQ1Y3lM6ST/SL74dc0EYU1OGDM6EkDaMS6TO/mjq9tVlnc6woaT5eHG
KKowPfNbV68/l1Rh9Uh1+xGkYBujQRQzmav0X9ZL4gnRwtkWk/j/Xp3PfPyM+G4tVjkD0SA0yVRU
WfZwLOlTa/sncTQmRBi/ZM+j0ZnG/HMcSN8djvO3NfHN39huhptRQj/dGaD+0ABWLyUUwP/eptiY
DA9QWJkcbHFJIGN1L1M5wPNvgHqOd27pbj+O3WpXFtf1cr8fp6Kjbva4MhM8ezRnt4ZqibcmWsCM
24hiwy2ujX3IE7RafV/AMCGrvxVPalxM391/lM3GHfRLrfNZuqM/P7jAjP/RBVtdyYuLQbRiSmmy
VZkWRTQ4AH39GvxpfMdlLHNujGzvQpiUOcnlUgqUQsKMDqJ/QJOqYyq0LmcIiMWM1CuykOmNYdSf
Fk7hwRWs3mYHIYrVITRKTBqeOdybFmgfq18/W+mgkkY+UhX6SGXSHwZzskQULBuvVzEYO05ES5MG
z6AHi53YmI5od8zfN8/g95pjqQLcglQbkBQ3yTaKLfUiUd3YdrIz//5fAe4KbU1pE0Kypy0VnGno
BfAoVBsPPbW5NuoiMgzroAnefCsREyffQJgN4b45PKkrim7rLSGN4CA5y+Xdx2uLZRVuaTmKb/oi
4DeIBx8QrlzKj8Jl6e2CZ5Ye/Nnc1BxwQhT1zOuGK2165GaY5Bl3PWjPbuhCbNpIRe6VAP1HFfVH
kyGtGTuKf1SHtkrCD6PMbYEQIF6Cegxj0JRIPz9ITGbmUH3oQM2si1Pr4gAL8X+dvrDhVwmq4Y6G
cdG+hZOe3pLMGh8TkXSgcfMVQtcTujnsHHFyvAj6IBw6Uw0fEHwAV90i1N6yqsq2IhROpblKeud4
y9rAUuio6HzPBhilZCwQTTbVqX6IBcjN0cuYguPQfgsaJlmTIQ9MWRx2yqgX25u4fpLw6WPIj05T
1vcjjJhnrBW18WaFDHj6TELkl7783CK5edsYZrrL0gBthTGMx/yr5zfmsGnMsHtDA5CHqcCE5nI8
Pxzlxoe9amnhIKvA7Djm17U0G8uic+wtX42ILVG8kmbkmiz6X1UogZ+Bjeq8FvYBlWDqLl51wr+E
I/oRmc6Rsv0BRLZg/orfTAFocpBhZMPKHcJoi2LBgAqiex9HTqZxYDAkgUOfAyqnIcAIKz5x4tEd
iwv6V4ZPjWnoBvWqyxNIBs6/vGbcId97tyzM3M9zCN6XPK9OkBtRzAiYIMkOGlroLqPaLfdhmCTI
UqQI7Em8hV8Tp0p4L2aTG+pbWzATF1/gA9vIt/qROyY6pXaxSzBGrlheQwGadkqdbZYW+J4ZdEmP
uv2nE8Yk1k0etHdxt/npJomMu3ArOPN2ZqoIVmkEMHqQYD4JI1+09R1JIC6djH2pTVX6rrOCxn+z
VRwQYRCch0oEEDejw3Menr/5EzbDvo/mTwYmcBHsetm22oxbOMJtDm3pFuL6cZTsRl5yfO8TCa8U
GYhCCdobuuoSaiy9WkeNH+fZyNW4XtWjOGipegd8G7dmiLNYjr6jNmOiNjCkbSB9xDl2JtaPfgec
bSo6vGCDjyxsHSEMcT0YAinlft4S+HMeiwCRs3vLMsHyHW1WTynuhO2YuYpgYzPTWn237PFWtWSr
C2bWOsejUZX2VBtpxWTkwdgHI9zW4S4z5E3l7SI8OkBsCe1tD4Z9uNxvqA14ternE/ntQpaju1i4
EkIze8bFMqPC5lFZIrMxOptIeDZLAEFyY3DOU8lyANVNVhL+oDqu9Xzcb4fdBEVlimruF0/tiyOI
oKtngnBUPiDEUbdePLJsa8MqHXJ4O6axJQEDEq44JydkkHU2S/2bekDXNeitIQFzaI9hQdUZKo6j
folKc9l9MkOSHrq1yMRwAEkIREq2m/29FPaimlg3/1PaH4yW9KtpOrwKVnWkTKwKOkuPI4kzBaMP
LKKBLORB7CKwa5T6Zfcv7mSG1HlWVJzznEuhl5yqxoKl0zK7stRIrZu5or4l8SJrcbJAskcUAnCF
e1SFNYZurE2mYB2CyLWwAwwNYJLZUfToJuOCGVZ7AxDFet5EdP0O5FRq8ezDqSUrsSvh2KZRbkHf
qbsgX5eUmHO9O1QM0aagJ1jVaU4fafTVZ9bM0IROOyU0o/fz2vtQOgzXkvybLApdpbhhJ2aRB675
bkJdVTL49LSxT9DbQMOup3SNy0OXendTFUlxq8h/VUCRfx8CeyQJj+OcGl5BIIYDcA6aTUQ/5F1Z
DruMDeWdqP3rxfSEYaOq6nCSpf5YITUNxfzMd3M1LpBWYN6X2I9CroQLaS7wiAkTCM63m/Wvh2mY
PsV6PWezJcgcd5LHnESjsKPzOqpGNLpJxFan4clEqAquZNrqOQEeT5EWAS/VQJTo7c+4uXc6nAC9
T4Vrijr8HlKm3DZAXS/vlOvbTg0sZJq2Fpcz9FyNzj/iey3qqa5NsRkLoDqWFhXTmRWwFGrsWdfo
hQ1Eaelja9knwq7XPpjiUVfu9WSOKcJtZUTtmso1cC+0bR+CodGo7w8CxV1bPPJteIkOq5TL7MGW
JIE1YfTQo3+Ymi7yYVGeIZ6PTxn5z4HFOUBndGLPq7QBiiRQyixSUjnaNU6gJCF2gQaA0iy5Ig5p
2FdDYdIqXy3U53ZbIlZJXrGY6kh16jczJv/JNAuHNj2BTDzV9m3jwtDqCLB4Z+7Lu2u2wiO33kRA
AaMwtYVVcOrDt0ec26wQbjtpq4JaEXf3bbJHGk+3eHgYDBD5HDd/WfTMnccFe7Ac6SCdnFyY4Y1q
Brys/2K8+jkemwQy7gBhp5HYfRaIYvb8PiASpDk9yxrz0ZydDFolPJ16I7qIVaYg+2NgtLYts0ai
AOAuvGghUVK4/TwbgufTs2hLuCi4ngK/uEKOMIi6N+OdTdyUv9XFckNRgz4QTaygusliv5rktRe6
yYg0IOHl2VL6t+abgn7P8PN2mHH15fbWa1ktbYbBggKOyQ1w27n5KTV1XNjft7/Bas7TlGi+xnQl
4oWipaAg6NhQyMQYCCB5NEGy3g5FQG4O5T+WMCGSVP1OT2En6vWWVq9ccw9vXTjINQiVJosMjPq5
kLEE3taK5gDtwb9s6AJD9VKRDWzFKUAh/yNzmT2uDSi3YsBf2HlY2udWW3pgCAsnwTlgr+gL8q95
F0h1QXPojQBX05jTSaM8h3Fjz0MDEVTsLc0J4d+LKI1QN2C1wxYbHbiRp1xzCWuLFJerhV4FRP5C
GIvFlxYwywiCgYYDGxuh9fxs3E/+rJhuuO/uoQMMc7IRgS0ssV11Q7MZ+Gr8cAoVQB9+Vqr0qHEh
HPxXKsKGYFdvuGXt2ol7MQ5e+gGE1BSeOXWfLcMBD3Ibq9nz6D7v3C/D2SXhDy38asPaVeUy5C4E
kAdVXebwScpUpKt+HvNlP7/1p8dUklzDYgK454ffG56QZGyuDLi5kajLmn4fgD3bqpDVfhRexVnU
Yv81l5rmAmYZcWMs1mSogaeG02/a4Flz2sPh/jpkXjhE5aIvmfF9Q5n6FsDKJBWaBh8z4EpnUF/6
M09kAHQwJAQkeF7vvlVM5qgVhbfaEATuM06KqjlL6YwMC+/Qva2oF/yoT5kg37SET1qzgpTh6B9a
TlWVpnIKOoUAhHoLd6OVXdG3MRXURdEXzW0C9QAGCJ/L00YJ8vH/L8tWVlAQpbCGT6ww7sr9STzL
5BA8alCivZHhYuaTfWuYm4KxraT1UBXiuMNcmeV2NoKydJDITlZmaLAmX3vhK480svDZNIPQvhg8
37DwhM6BZRJE/MzpjbvfndygxGmRPruNYqdJX7M1sLy1V1/TKZshpCekMTD1daFKEJcUw2p9/Na0
/g0C3aIrke1swAP01iEPW2gtzHE57Zz7ji1T9Sr04Foo6spUWYvywrcLV3tyHDy2z1dp7Ex4IZjc
B4XwOG9xU3YXB+plcAeMqt4/76QcwICi8hUyY5EAsGPNMFDtvlWZg5N5Z17viuadKD0nmarTBntI
QnWaQMK+XXqeVFcRqjEyRtcOQ/607Xt0IsxgOvWnxRC3iaw0S81LepIWGuCi290zebsRFry9xJfo
gZRjOrBajy+9I+93bdVhuTM7s47YOU9WcdedD220cYbnpCLOxc0MtuF6T1bYpQadn7s3g9+kNePz
tb1dt1wlipbCzt7rVSkpb6NO8x/qGqa3BI5cP71+vQ/HxLj9LWk7b6VJUTil/zvQMcqwjTyCioSp
UPzu6Mvh9i8DW97yMC54l/tmyjuQTv5QjsT/eo41xUXtjANw9YGykxBd/N1aP38QD0xcukWLqEP3
0yaoQE3SR9gYos2DgOdAPACM4mTa/MG6vULk+KAOxDnRe8EH13l7q0vbeBfDts1/eJRsfFNLalsr
49J18sssTqrmAujVtQ6VZiURojyhFkEn/UQ0xwbJWayvE+HOk4Y4+hp9BhvLVIb4J+x07H2SoVcJ
S579oxPIgQgXmQBqTKSNQqmX03qOezVAO5XB+jDrIlxeGzLHMvf2rOryIjc7goL8QzRApsadIt7j
5UNXZZeSRac+4dK9GlUKlsKB1F4QLMudHhGjzjv96xMI5Q5SiTGcqP/HPKql+rpABx1SfcaAcJph
acEcN06svTWdAp6E+hxYMZJkoAbmBdVmtfEiOCEvlPpRVhUuBhRkYysyDd8b1U4H8kz22eWOIj3d
g6mdJUgBp5dZfZ0Ld6ifdgarWuksenqVneVCWWa6XHZ7N+720Qk0BUZBEr1EJaiydiOIZguzsL5+
6tlkpihAswz9tN5qZWSdOGliY67IHbE5KWTBoUIdN1h4p6NGp2SRFO4iPHDkSob8GbXNceumgmv4
jUlDY/bqL28puE2VKa9nTiJ5Fjh2R0aQAeGQ3CmOlR+DgAWpMh2b43xyWj7Kls1v27BQh68m4m1s
/66VkHJ7Xm6WcXi3muoeu1mcaN1fmTEXgPgel5/0HubqT4JyftsY7rcyqBSwZUOz+SdAVfzT2zGF
Z1TYNdgshOKI/3nVNgc/s4tjZ/6RFkedSQAmdN45gRmDxOxcFauBlSO8xYYUDSwPCVue6akn/3L6
uH7BDhP8H2dYnTt/Pdsuvs1YotAja5604L8irD44KKGbksBZQvJImdtjfWxfG6Wm1EwlqXXk6bpJ
eUF3fNIlnztyOsYpgxRDtpU5iDPL2lHSL/AxWtAWQEDdBrDXDHysMqAT/gsRfXImbo63jlD4MKdL
58RfekHCW3fRhl0p82SESkZo+UlpyFvG6jbrXZPE4aSYL7aNQyl6tb/sTC5328itkEN6HGcsUB4A
DalFBdpSY9J9gk9bnYy5k1Jy+HBLoT/zGAMsEPlh9JBxZErXJW7hhn5EO/2Hzvv3FIEHvQZhkgUi
zMa7cKcXVjX0amQuK7VdoEE7aTFpXhH8hyn7/aU5qOPVGH+DE17PBX0VQoFelA8+qDrp9jfIjjoY
RWAyFPDaUrkcJG8IpnFuXc6ny+lekM4E51QU++dKEk3sk83/gbNYoVp5QXT+w/kU/3i2LJ1cGWAv
1D5FgY/uPWI0+xzR96XKwkAmeOuVEy/8vOJ6FebkHFDUmWEX5iDcsPTQCL+M5CZtFCT165GZb3GW
fK2qtqe1FR6JjZNSZAcNIY7xuua5JPV74BjBhRSqmseAsfdgpJqTEhz6w0RzZ7kYKKt5fJmuOBh+
85uQ+fNa70hIE9TfJHcCyIG438tv0czbAQUffkEBQ0tz5zYBPZvnp3P8OdtrZ1WbKjQvPfSCvJjl
ZOXUztLOKdgea3mJN7MaMCOSL5FCrx2vuYayACTuE6JnEj2W2N6PDvBAyPG2RQZxRQYGjHOC9LJr
1YamCjTfIvP81OK35iN7i+96yRJSGpXC51GImZjK2+LIP2BOpYwRA09ZQzXys9RT2BB5nuqhMv1v
GAiE7GrSo2xkiTpbffbj6gymswizwDKJA6b+BiRgjhjeWrKc2gZhDj6VOb4kRUg/XYudXtdnFfEV
WE9+QyAT813pgZjZWj2ZuzYK6VavnKk5joP+0TAmNqvwFiB4kagn+xCWIaWxxltSYO+2rmd4WEhx
DEFNo8Se60B05SV2q4z8070uOvUZzcbktTj3C1bnd3resYYzRJ2zA1n0wmFMfNNLDHTqYPSQTuhH
jhugE+ARcjvUV8lvZIqMd5+dl13+LmHOs7h2aU1hUb3Xc0UBnW6Uzc3pUIxCYRx09f85vSFoKfZD
bQuZJP64bR+trEUV9o9TgFrYLahD8lPUvnC5UhShdChGB8Gfmfiup8qYz6l4KNgN0HTcc9yFebyc
JhW3aFFY3SFXr9eCZXmyVPjwXMgFli0se1nQWhPij3HOjdUF0KzN3myO7wLZoCojnSKiMyRx+8vA
JZGDEzfyuSbhqk9ZnWBQWKx5WDcjrOi1Oom/fs35sk2Lhp2B3MzcSQ0PXcgZih2i31Z24QRuiOv9
QXs475+Wd30l4pwqqaHWEkP6wU4MZ118kBLj0J8KfLQeAYh+VRvoHaJKEX73u69H0SxHW4VY6Lh0
9GBfSraVMROZCUqsRBLC5NPkK+gorNZCJdUrKv2ueBs9YXCqH9RVt8cemIZKcbpM+nm0k4q70ig4
UdWeWYd9F/4ScYiX6VCyJ5/9FtuvCsODnNQxW6n7jWgdHNCLyBB5FqG10S3UJwstQ+ZMXTe3kjAI
4cfWe3tmKpkXidWDZHvi/v0LwZk84ClApSYjqlJ/z6fixEQru0EiBp5kDrcOfZdx9Abwv2N4nKn0
1jkSIyTETBN+USctF0m6eYjcxuNQdBxgFbIIGgiiNXVJ4dTbOqO1pX5Kpkrl7M10CgQvH9l1u7AR
Yapne0rwPSv79P6PNxIlwmZrjFbruzFicfvPdBwprEb2/01SqIHxpHSDCZBA0sVj1K/GYKEZkyPI
jWypCRkbDfhm2UqtVP6dShirJ/c6PRIrA4uDNajyCOAy6f2ajI+FPlS4XiXUomx7nmxyXWBkmjnY
E5urCTW9NolbcFJGncN0YUVjKCpATlY/6l0lvGeN3+zBuB+84/X8G2md25OFO8+8igzt4flFiPYJ
T+DlVz0nmi2Pi0cRIpPSVBp7bkaKH+yvnCubPZH3WcQcg4OfuicdUIZGmdPE0adyQjuICEzbR1O1
WnPbGslR9T1NaTm+MWaklJQo5wVAAGZQqsGGGb3LNnQ5RuM8gFoJpQGloUb2mcrW7td9ax9U059A
GFEbS6IxiEK7vjBMMZPl9r9Yzcga46MxGIInMY2raN5nSQnBV7GdM2Mg9FLuS4pj2EpgkdyQARWh
ndRDmAxGn/THFzoP386YcRVIeJsazML5X8UTec19LrGiQQymUlNV7DfPJLYwORmCpmP6eDvjcpul
rwe5mKZDqIHkHaLJIURorIBC9DdwIZ0y0tYAFoKxK/Iw5TSgn5YqX5cxAlsCNnYjt6r8uWAecDrj
XLpWe19KZgo+H1kpun4d5jDK9TrJ5mdbnbKnbX4cX+TyJUHAy5lH/d1Xyqkk3rD3unqfVjrv3Riv
oT2grJ5FA3J/YS04QUHypmOB3/YEdbFXbBEm2IdLpq2WnrkKjhKrmSzEQLge9tWs3MrGcFUsKMao
+ZwqeH5MCXdcv2zZnAuXZHLrbjrBNnWXJCiuVvXPTU0S6nScLHy9VQUMP8+5OchHHa7G61evQ6Wj
hbcBSHT5CMQ5ss/rEL6ZpaMchkOYlmSd8gPiDpuPKNjfbJmFNuNbE28A/v+lX47+wcC1ohdcdE6P
r2c5e5y00JF+4OIVHainRwoQ3VYVJRNqEYvpUhY0JdVGz4HN80oDicipiudH63/kHr6OwmnKrBRz
9GcqZejYfDEoFUxYVSuSnbVBPWtj1pm8ja1xwzpqDr1Vc53QiK9QOLSPCh+hMC2OPcdqPwtRaWw8
TlQNWc6d18GLb83kF96qg0UeR1aCzDO1rXVZz818ptTUhz8ZEE8rKKsw9k1Y7PNi7zHk2NAo0rIU
YA7rFyxJeinCec0IrWqQ1jlX+QhzWqnDcXr1jLSXF+N4JEhiqrkeDuSZJ2oLjnmJHoT4tGIBnYDI
S0Xo449DP2sa4/jmAZGOELrzmnTzQgucC+7R4uqzEL5Zcd6Lse89+/Oqi/LGn+eK44tNFgEgPvcC
WjFg8aYk7/Ev857W/0lcJPqBvcrkfzhqhyppep3cuXShRO4FvIfxarIm91EGQnI9q3q/Xm2PTRnC
TYKzy1Vy7aMOOuRfruDhEnPYtTF8PzDc/O5IeFtr/kXYe4PoGSYvD46MaLx4ZhNiKl4tbEDbj0t5
b9rQ4Dd2TizWQYM4Sz3FR7MrezCeP+1nlDNznnzl4BCDPS9wPtV5hQPLBuIGYVwByQGLIrP44E5i
V2RAjHFoEvCUXPAp1kor0Sz9VptuiHTKVdwxvtidwfnQt/p2O3ZxBows6X1XQdo4eBLT4fiUAgHQ
a2jgkQUtorY5ianIZkXXPcZN3H8pA5nSoHNmywIYKG8jNL3DP18qKmD5xpHxp6B/IP1y+trRnyNT
RMdHaIGO1YhSzSCce1yRsE4umYBEO2bw2UD0V1y5OafSxp1yniMXTBPQxhMSk8oyWwQCbib+Y1Yb
XAr/xHnVDVvMh4a5wCPEjWdr7ViNQ0T2FD11e1vPJG8U7JYnKhJF3kyB0KRoqLeKsSsyRHl/Je7O
+WJHMRP9gkybuH/9MHMDDD/HT8OLOLnPu2v93o/0K99L7U93ZhiBlQDXSFy07Y3oW+CTkzpydRQk
tkFGQgdH+KsRJTD8/xodvW3jrrSW6Y1fF++6kS3ixFIdqX9SN3Cl1fGp/6dbpmemJXkAKdZ7Ab8f
IkqtOcm0nJZeKyTPk8vipGETZ8zyBe4biKix6JMQV7TWdNUObWVoHG0avWMOcH9nA6JcRHd2haRE
YLWAXeVyL201nAe/h1YJoUWuIl8PDj/di9fOHeRiWrdZwljKrl3Hrwak7MSVmOAERO8dhUCPg8vn
omf682l0Msry9ed7wud4QehIzjAmBen8/SVHMGGzN3a9bSFvHHD7wqPrjUlmBfwtEamEKjwqIKqB
Nv+yAiFeYoDB/92FC0CDTzz3QdNjyjqjNxZqjr9rHHnfQVwqHyLocb5C6UAt1C4+/2fQQsFZ5hru
mC69gy5Yv3nmaPAkcYJsMzA0lqk+rhxV8/HNR+sKJgj/pGtrYsdcwtrUL0tGLD2H5hKNeXaVxhjH
k+aZgfSISCXIRK0IbDfc5CIX6Cdrfcr87DebF+mYLorI95DblvesPVPg/nXI5UEm2bLmwWgsSc2u
2NcRwptWwXWM+9tndOE94Kc4M4r2jx3pM0EstoR2NMekSGHoSMi/WLXq5asSuYdF/ZrduHpqHV88
yz8PWr20qLoTWWClaFzHIzWqQt+4xj1y1b6XN0hT7UwMyzDaYVYZBzXaN2szVeLwuTD2+AxIPL1Y
HQ141DZ7sXyK1VfDOzkLYN55CmdOiVThJdadYRzWIr3alacrO49WCFav0dk/6+pix5gZE2qjU70S
gXZFb0UWaFsaWxxVIwlFTOIYy0WvVhFlH1zDdq518c7BGQZyAy/kN9DpCYv1QWCFIiylOK7FjMXY
o64obaWYSoROu5Md1nvGJqu5gxOSaiVOkYCTTREjMzzMtctPR5XMkTap2jV8CejegGCKCcG6Qge/
xYaE8IPCkf5mz55PSUgI+gvDK2mPO5K8wTkD1MFsDxW74gT1+qW+4owDAC3obQalD7KZZ+olMb1z
1eZj1jSsMao2iDZIbS6jnVPlERzCYp6sJ9gp6KaZ5z/d7ncPji1rhG4xLp4Xk16BFDmgIVA1wl+T
bupff57aq0G5dfB18LuPUhtm8GlyUMMo4WJTf5tKF8kFeJnaEXKkXZpX4xRJ4sbF+BcUPe6l/8hD
SdA0plgLzZJ85M4dMh0Pr6zJnhECdG9SdT6xsXYzMBOGw+zXDWO55Gt1fFfP6ODz8au/suUl2Nx1
DKPZ5Ud+B/NVHaeTN6yHrWfR9ygufqvviNuCgLzsrQzvwC6wJJ2nWqFTKdHPSYuxR+itI5yDKW+b
gLhcmGQQU1V/AjLYxhHjE1c3Jiff2OI9goiGjJ8WWuVbE/xh+5MP9m+nGWN7ymyX9x4CpKs9oLRX
nsZ4jb4v1KOuzpGuavIOlvLYf+B+xWPAw9rYkTxpOEQvSdEuKB7MJmuesuu6sf6tgacUkGRJ1MXY
muFncykX9R1VquIgSlTtbBPDMV3hHggx0iGIZJMdsAxpsolvjfvBm/orxC/Oil1Riq55MlCtIcEc
n4lBBhEYRbZPhQm0j6kYXc2peCabEjMhTTiLPV19m3quF6akeVrn/B3A4Y1Cyzc5fKu2Sa2FiCWL
1i238gIb/JESEIh+g/lB1sHl+dhHRkiCOJxs0rf797OsXm9HLI33YrgZtSD9ngrUl9+wfklFs/IE
4bLkNS+lDudsCpdEDgtivezMz88bjYdKwONj57D/Hi4K1s+AxPbYe0pWJ1Oh1fvkFtFEX7a1XNsN
NFXT3J1JdZI31EQkz7jpyYH2kt7x/Gd0wgqpqmz6mihyXpHPAP5i2ycVTl6IdgT15KFKQzDcPjY1
hCg1vhSUTUSHOs2lLjpegSiQp2wC2I4p1oqaGEq8WxB6FHa78TcXXyV97mQlp8NmI1ruTXSq1yXB
XJeY9Fh9jYZueRH+0ibUuQ4x4m7v8ReXOrUvv3tc9GitkhOKtxfMlnZxEi06i0mNtI49cCq36f1c
vxIkYf0HCcWwinZD774MztvRg43FZIHbhMu2EHbonNv3AUTq23FXlG0t3SkCCcN8U32GUXgdMiKT
67lU8MxytxREAR7W6dKRVd217NgQrvhuzZbPx+8KtmvvtPT7WHEfFePFQ+TyO+pCouRvJ/2Z+8hK
qokE2i0DMpwyBsm+N0i+F0WQh4945KLwXmmqK7hnbu/ehYQK4RyJSy4sw4AwGAog4nCJK3KNxVyX
xm0GVWqgYGQPaP372gai+Jc6F/cE8TkOcHoG08dG85wEmc2u61vf457I2jV7MbP/bmRtFJm1gBAT
l5SF6sGL1H7xBO286KuOrXV2cUyKBin37vq0PZP3g1U4DNGIPmrXUHcieZGvW4hyDK+z1EZHB3kB
ByGAu/UUIq8PmUWIPTHQCdOE6VqZSp9TYrUjjIIH1tMW65iWLImBa+rTWNgca04IIoX4Lg6CqpPB
vfeBFgJAwiQw3TDDAZuFPelnZurq+fozDHw4H3L8ISs8mZcXf9V2lQRJ0UuizqdlE7caPN1epmwe
WJf1hO5IyCxNTVDh5FpLZzCezAOX2akb+d3qUwt7zRCaLmcmmxwHr7b7oq3Bvdfil3CmBFYqI91n
HTYr9tx9yjuY67DjOY0VmfpH0QYbOeoG6TdprTQImBkK42V7tjGyWjdg8LHzsZZ16pmDPYG7X7jZ
wotEx2rYAMgHoRB2y6jMUOysKkH7qtiCgM0zMpI2OeZFDS3bFzLeBGp3Aefuc4AVoFB0z4ZJczpY
oaF+eoB142Qh0UWZx/GCMrcTF+RtRIHmZcKRFYOU/Em6CBzDBEA68m5KRyFRgjFsPwOe2FsB82by
tUF3ZtbQwyVa+mLwu2jlrjDcpVsMg/bItJyPmJWnfEyUaUtDJDO6hyz+Mb2omWwodJsaCAA8r6GE
0J7M/PIaVnclvnkn3lcxfCNAFclSAdjK1QRupmAT8tZSoMyMv/dDDRvXOFADX1T7yAVD0RT4jGP9
QcAqqUnAU8Vrx7oTuoh0PGJI/fsfYGTQkfwqZXBfNBuT6mrjZgCMCGb+EA/8eE/ZJnIXginW2lz9
jmbuBMiUvRVJZlO6Z7WsEI/24ACvp41EucW4jzw3x082JO4CjPK25k1MYCKIW08BhMiibglDXDY3
/SRUmbhuJK5pGCEanHlOcjTYmAHQ62axFazo2H4Tb4wPJ3NUxG9162qjkSv6vgVwpH2BcfQeftvW
tQsmGDAViCgsY+Sxi/Kfkx8UI9hx1pHqtqhL0oAKyUzOpDR5xymc5kzF1WzLVhOSsmfG+nEliTWe
+38x4SmT+1IbIbTbHx6HTvSTS9naCJpIeYfo3GzODNcx0+qSkchZt6p+nTR9qfbNpIPDHN0NrjqS
KzEqAJLOzrex4ibRpeiaGzH4R42JHh0nRLzr/DVjcihX0i4nMkTgk1FTgdmKTYxxSs0rDtNXe03b
1GOSxm+MWWcEU5aIVvZQA8Js1t3A9k1UE0+/tY5TWr4lT0RaB84kl83vlIvypWncRgQE4yEYvjFo
tud+b39NhxlF4nYogl0DEFt2hLgx1eAG5n5+VQ/v8pYpL0g+b2E0CjGkIGZV48kqpkknv15aTkwI
vlf7cHa5V20haNX/dKgW6i6RHHuZaVG6hWvaFJos24rDfCvU8+ASwwZp5fpXp+xBGv4UNH8b0cWS
FY17CI005sQ/e+jmNheRet+/dnJioB85JfhtkwuFV0SlRzYxXSf+59Hmw0hT/+MoU7VxKPGfjjxy
2eihCLbSlA4nVl+C0m9jZpZSrTYs7IlgwLQ+tjlFIhi9YaqwdaIX6ic9+6u4PI7IxGkNBkm18Ctv
qgliGKksgR4cHi8PDgW8dylFeM76JT1FeRjbt/n+u2/Cc81st9AwHJYIKOd0VMmbALkKWfaXodZC
UdKmGtsZbjl+INb3/CDq6kMIJYF7vf3brPBmQhHs3/Y4QSPrkoVmIfuYTSkVbm/7TzRKe8LnELEp
sG2Waf8a9TZToSSyOKFCAcTEmoOQvi+QegwG6+Anbp5Lr29ks7KOhZZHCusH2PuM6woQi7j40fS4
T4PkwzeQXzh8hJ0JhyHQs9+xC2tjhXgMxuR8tu1sIGb+XebWWM7sA2oCSVoVWSDNlYCNdxMuhzMg
tikrCstrCGsxRmeipDwNsq7pDY4NuPuYlvOK/auT2/jOrOEOTLDpiRgCkPw32j7+Zyo4ZVO0U46E
XP59TqeVWN0xXFlRHpNrbeBT5NZwRfrWkcX1NpDQiNYApZLbsPmRguXry8MHHqkkYqqjGg83lAZx
zXtIpIse6c+RfbEXSGM7vhR55Rh4A01OOvU9FRN99WRP5D4uk7t0WRiDHRU8mOCM/YQNFyRmdt9R
kDVeEN5R84Yfxmh6iYv6eFq1vNabO68GiHcNZcyf3sX3w0kqrE3i9ZKAnAzVamnbIWQYlkkHziwB
/ZINDGoKSc9BrblHx7oISzywZs4Tq/liseuEl5z51SGFBiacqMhikEZiKfuBVmdb7aA7PjGcbEG0
xlU8pJA3/CHIj4xf4HBnCt9HYm7ckliDqKORxBYOsIqzF1A4+NL6wD24hC6qOa2kQOs7YNPad4hx
8LaGsUKlwJKCiDfB1IKNk/jyi4dXqm23nKbU916B7kfSUXPFEMeFicHXXNKpSDpQQJkxToUbB+1F
CvHOqe3UuHx1i1lNUpIv3UZydlC/q84rha/AxIgoZEYA2VyZ7xaskggRbBgm99qu+8AhmyHYvaIe
qK/xQR1GpKKozcKKoSBsPXvu22BQxLWFJnCYukzVeVFvRXzPhdDtxdO2aCFNt9uMW1U9b9qv/UDx
+oHiY/x8f0hwYXJFSVwi3q3x4syPZo66Zm05uiaDBGtkZBiVh+eNnsGtR+9DYTm6S6SGeFUkkHjq
BAu1/rAxH5+0C6DH1Dmcc+LQ/mdqqoPARgFGFqQud4CZkjw181hjaTD9DBWaVFnzSgxwEuLhozZI
pzs6nGMqpfaPegx4tFVkaPZrnGxLAKdI6AlP5xfdIHTgac+nhJ9O5Wf9leA/HygIPA8cydkhLaad
KOyRUU5SDESK3RMUp5YifgBg0CaL3KxHZCLP7pgarX4JqBQDJgzf6/tPgkQ1nWKpeT4muz/KYX1S
fZDWcLacMz5imFXK85wx7IV7otmVVngROH+D0MJYJASvEKHJZN9djy4uf/YQn7OnhzOJJeUZAH7i
mrrS9lm330E8MrFpvXcifvbDATvy51D1Ibj1k+8mTvlPjm/hW394oxB+SwFtSC3Ft4ix4ZWhM2cr
HASHycJJ3CqBzGTx9fMYUZ1hcwr6jg9JoY7n/kBYXWAHeABh5vzqrfT3QVJmiE9sFnwHvFHQhbx9
nX1eoiLzFt/aOe3/5xzQMbjz0csXAHVPTolUOB7uE/qAQ3kuZKEcqzzwDHxN8Y5LALBbmThTyRBt
+zrjfevxkVI4rgDpz79/MewvGeZH2E3CzyDCU/8zSG0w41w7T5bdngAhBIzqlkmnynaxnDvgHeYb
3O86ibtRbCpJELS17TbJey1Y5sZ06fqT83L4vHBcsiXY0T2zTGsdz5GSCKTFGLHW/UVz0ujWZjct
h9FATEvRzrjPmlcoCAn5fVqjWH2Zq2wIfGXjOmgDd5grkuXbSlGc01iQIDsboDjO/FFRmMuKs0qt
75AsY0USAHbw4zo8m5R4gEc+wHonDWGJmcTu/xa+wKka8mptP14aUhjQ3fA6O6ka1VaRQ7lHxG9H
yUCkmpo2z+Uxl5hsKrU2YkwqAYsfif4ojMJ3R/6+r8KRSzlvcVsX0oRgNsJIqNZEypde7AwuqDUn
f8TLSLnkJHANoE3B1IVBh//IPkgN1le7n42l69yUMfsKgxp156WTXaeWgSrT9AGUlqwLGl0MqgSq
2mwYU2eCW1qPIQuczLYZHuewJE+WQAf5QbLju6qff537rjwlBgNEfOvJWDQ5sAyvfd1UYObV67ux
S1uydesMrmNisFX7f6/cbGswtaL/iKGW8u3yi4+9VcCW7qVpLSCAIcakQ26l8DuaxkZ90ev7CNIX
W/dHQ3SnUoPLIdyFOi4xwKudasOIUo0EXWLNVaeS2H5gLk5vdbwMXSl/Wdnwo57xeQ8B/ReG1qGQ
JsUAtrBQU8vDsRX7QnVIsYmS48rtnlPdMfOfv9tB1z3dumPZB7gzdszlqBS+cQLjI78bDM+MYJVC
7rxqoN76Bpu8W+IsH47Vx4G+FpSIxfrVrno/+ApI/O7zu2ViM1bgLJZjBt8Zo6hYKSYdkIDxJMAl
iAHaH28MGySy7s6afVbPTHSayB10tQsXu+QI8sEg4bHe1SfRRrATTCSR0kA5gi+EUdVCpVEn2HDs
jOHon1giZSNWRsvayE/+1hKffmX8QqEZBCtE9l/F/fkuQLu36XRoG+575de8Y0u4GRk67xZP/Bwm
x2XYf1//ZRT5H4GdLnzCSUBclC9TApcH9mCQJkruwMqueWcIJ42p4lRRjRpDYc+0NVVRvYGenB3e
t0pgQZMXPcML/AYLiqWQ4G10WmjvWowP7hlVzvi0O8LDIq9NHtyuxwqQpbjBueBVYOzd4S4UY0Ap
Vmr6trxdsCMOeev/nKbD2LG/83bWfSq8TZtrc3xZIFnnzlSQ0XdVbnhI+vIu4L/z0IeOYYZWsTbP
re582eQ+UDnIr3lVP33tYDa+JL9+9NtOkRCWdgg8LeKcope8i4Ak+C4cxZG4U2eWftP1Xhd21hL8
QD+h1T83AQaGuI6y28I/Ay/8W9bkbHvgjNc4Njabne/IJRAbVrnNADB6Lr8eBGjnYSSWfA7PNEs/
wH/FZUEOUfEwITMVYrZ3RupcLr+7KsN64R2Rb3rpoaD2qhAh2I40NZ09XLk1wuSWNxoos727762l
RRmDtrzd89ftsHM+8Gw1R7FEF1EKQtIfQilPVBQyouW+2K5a77rOsPs2JhBkOadZ4nVG58Gzx/pi
LxNyfNpRNbw6qsNLIY/FR0Buw7YqSAue1FJ6F2EWiMSLl0h/6v9BZlE4dp5VkT98JLcQSiQ1BHng
a05sWT6jebEDnMUG280wkTsFIlKB0u4gKaAOeKlxD7LVGe3wcnnfdgv5lOgXVnkcu/unGVJcXYa2
Vy7qrbxaGqOv0EOJxwyox6sSWrHqyI14mPwJY59a34syADVhzT2fzQJQtu/7TKtNpVvqZqyR5FgL
uSOnMVPM275S24E7+cwJ8LdcTtMlYrvuvQ1XNAh2k8ZvCqJYPJqiR8wdvEoK3VCSyetFIv5ZdfKb
K7zM/HRN74X/6sgNHr4SZy7Sc7InBKbmtH9++0LlL0js7/xJ1eaKBs4bOTMNGliuUC8/ztz6/5PZ
T3SjovGFN7rjxT1F2cJU9C0EfKKcCvz9/63+3gORdOIoUUrm1Ks7lFdoOyzTqnQ7QowZJGd9SSVY
bPLa4vsUJxH26HYhkvql/j5D7l3KLB44SqYPrwQx6ryg2Tcp6m48LdD+nwEVOU9fWfwNxMdy0xXi
XpCwm6wRfyrmWIF5U+/JB47mGtut0NT+WWVwCNCrb7WTZdSAHAybc7Hvff5k5q0Vmwx7CAt/FyXD
tOj2bThAL1BjReHcMtkQqvQJRPkHSMpvIv4FqsGYMhSF0QXSmyq2+CmBnBvBX2Ng7nBLNjvOHEWT
iXwI0Oqv161+xUlE02AkOByHrYVJoonbltSThiZ5wwnqsg9mfRKHhdF4Ry5UvbTIhe4zVnyRUxRo
9dH49zPvqTwUBNLkw2imedFFV3euIRyY8NR247pV5A5DTGTXXqIUnCx0TL5GJigMFXgpoqx2TtRW
6mZ7cQiL4n3DK9feiSpOkmasTon5YZVPAvRrFJ7kfJE8OYVBFUNxRdzkL0Mabih7cCOG4ciK81k+
HOj4ScHx/JvoqlJ/5783WYlVFSfc1Vvgu489TXRwzv79H7L8e4ne9GP613trpwsn3/Yf83v/TsWW
9UTREWz/X2XXMSEpNhABTGCIvZe0qu3jAOFyL/RW9S1YMPi1OdX1ZQaUOhKTn2GcqrrknllGTQJ6
2Eah3b4bAGHLJF2XnszrsDYLtXpENP5FNm8TPzGgsL9dEJw0ks+BfUWcCYXUeIjojSvdB2x7sqjb
mhXaslzRj/FESlrNGastD876qmtfeOAJUp+qsXwd92noo9YdNcOKyJhOJFPxid2XAlWk4KKQf8jC
E8zZ5RVGzPpZQ4FP7rg9mA7NF4tBiu4kpAweUoookwO89v2o4YcItbuMBwxmFJf6uvyz/6Slwh7d
uimO4T+asbMkDSQz8WU61g6JVU0Ljv5ymIWjf4IgOHpJ9yUyGlFb6X/w3CaK7IfLYdSoJ8pN+h0D
eduPaTOqul9NF5W0PIy1ikgrWucNKn+cEV7bcYsEEoYMhlXq67uCZIeF8Q76Q/qqcYYEIg4tZ5bw
rl7bl2SAr43/iyvdoHbwK4pUOW8DpY0Y0E2mgRT0v9NyOP1V30KSsnJFVSHuBclM+BLxp5FA3uTX
Hjb+ncU8xs2n5Sngdt40uuRoeat0hfejPxYdMQYsvNPj0aPzfMPnpthwnK/qlo9UWK1Igy29pKke
rHJ6q5d8Nb5UVbYcgZlxnBpPzrxjNVmbZ5qCo5WBjaQmT78SLJQNXAnMEwR7AQ9D0UVtLiT9PZxD
3OkZba1rYKFmRgKy1ZRDbvaf+w5Ss0xBKthwJTv/SswHDtvlTziM6s0BkdLBwoif4Wup1+Wn4720
dMOFCjy5FzrnvySQTYKfRxu5noi6oVayKAqUIHHfJM76xN/A3jAq2aQv7j4FeY295rHt0pMl61F8
kjkHMzewFJyknv7I0QccNn7DYEkh8UkHfDvAmeAMDLXaPkNUcFWuUj4Vu9UoaVbme0JFBA86AK0h
969evw5jm2aYAuUrsAe6lGkiyATHtii0U6WaqCQLTK+uv+UgE9Yxy6lK0tiVLr2HwmPPP8/B1aRB
oUVOhGTKIblGgahNxoK8S1iA7YV1Do+oS4i68bxVh1tevYlnllm9pBJDbVpjC7hGE8g0hxAP0QM9
AVVDxswrxfithxrU+Lnzwf+ttrW7P43wjYQIfFXTj3yXlgbQexOC4rBpyu1tbOTHo/t5T/t7EsV/
SI2l5vYDFIIy/b1OgUz+mfj35IDpgSCTBPCVD9OVcWPnlHPyAtovuZZ38FmjGnZVcLSZBXo6gKqo
RM6CXsCD81SC2T6NJ5EklnQ4xkbbwVrjv6guBTnuMydwgjz3UPcT0a52CEmz8rfitMNgnMzAFkjA
ID71zUUk5D0uEN0mGNY47tE6NaOZ6xHRLBnydBDgtSXOnT2g4m7LP0J3HmNcmjBN77rtnVF1Z8Gp
xgQNGFGwojA6UMdW6QoIT4W6wKSg/n4VPIyC+kQ6+Gu2YRlbfMAh/xXiw6V4zqg9B20kP8v01FJ/
QqJ+1C/bGIV2wBeEN2QJxXNRIO+4ZEA33woHbA4xzvPsZYLgj1PFd36sl6FbuV4PBIlgKHykzy5I
zOpgPrHzFVGi99U1GaaC3+9aYFrVnKhEiaYAWv5vZw0hoc2Z/33ZFnTDtB/JxLzcXZjT57PsdDot
v0aLgPc2y9HgLqSvWERo1ixTQNt7y486BASCpqvnItRGAz7UY/sp4t2/pdudXWJAEazr6veE3uxy
nDtVoX3RBNt0twcWt0/h7UgkSZjYTAkKyUHSQuxqV//sz7pzaVZNPzb/CLVyQpyOfEfzKSMqvX/r
QHHmczT0qk6gYS+d4Sjvo2rIB1Xr4vu4RW9UR2KnpCcVZMbGOlyRmGhi97KETOfdGxfH0xDq7C+b
CvqN0BOpO9m0Yhd4OZfmHqGSK//zJKa3oTrPs2bN+YiHJpTsTtRPTkX2OUF2Z4O8bDwUwUIIUHIM
h/Rhd2/E9EUBnVYBoHIXnfsh64Z80wffWkuLJDtFKj8SxHpalXoxiuQYaxBG/zk62VClaSispuew
A4CT/K7XqHQ5OPu5Pm//HOoFzE7mQH9aAK9OjQUrNbeZsJtFHPky9e3yebujFR+2KV3p7TOiajuE
m1dLO8t08FbXBtLO3ifoLCgOttCkz7pdH/NxEnlDEDoSYj84nDBCrd/yNfSMHSEKm6fdc0wTwA6T
OIgAquaoQgCy77e7j2gMn4cfEhggb4uxj2aegy2u9Bl7MuHpRVNXVTbG20CxkPBqXYdBJO1Vk2Yc
oJkQGN82hNSAeNh+w+NTtGr834yp9Nm6MhgKUezBpPaWvYWFK+qBSUL2GWRk3Dlrfx7fnS796JTm
vvINVAXxrE0M2vPvEJhqP7gtjJlLA0QnlBIuN+GWk6TY3jsceAXvYdrqlRr86H1qk8H30tGdX9MU
mHattPV4iD5EoSrOagCs9ZlDfh/3yp/O737p2gTNwQfmfuwV8tsXTrF29438cc6pyHuzltrf6Usx
nLIOcHlzT7PFLzFEd+C3WSanjGkl5BBOG5EVMfEowHeVCJhu2Dj14tw6QHfURaKLmarrojRREWXz
rs4kkvfVDFb+h4bKg5zp3oHPZ8ggefH8LSQSllrtxhTR35KBb9FQ4G0p2NciR0Rv9XHNfP8ZsZaj
jHwXJfeH0MDa2VetqbptQAiTxq703e/y/CPjM4oGuv7xxHXZaP0RGiyPoqx+mcaUrT9IGw1Zgqqv
VPn4lzU5FELaUeBWBQlKoxJ/P/2cDgAr9TzqkIZYm+uA4k4GaBk2braptVL74ykQIhQi6Q3z9E96
t70+JgqtiAWdJ/In4r2JEXIzllmmLu09hK9B0/a6Wsa4ZWX4RKgLM7R3LjhopFpcacKcYNg7swnv
v5EPAwWkc/gNLbxMpOECBIiW/Hy8QVivqBsrBuaJ/d3jL9ylHIhfO2KYM4enYGyubzUZ/unSI1Z7
Baf/tqg+mvTBADwKNvy3dV33NdEEyflJ/i1vfJcYn/ZWhTvqXS4pLWv6EGuugM8uwW+b1JTZlmif
CryQz5OBHOkxkvAe7TnO0ZfLemZ7k2nVZRM3gGE+dvsIo/x8ctsZg0yTgpTkLaoNGHjT4xmCzILK
qjsGfQMTSAJR30IK/hT+uAIvcvWsAOSUl6BfRGOxbHY9uq7K1h7TvlIwzSl7uSR35K/3mRXnevpB
2fwBFOCb2lqltQr/nCxT26NAktJHtuulHfsrINaODZcg3K2+n4ou5wEIBA1FSBimBYcTzMci4DGF
2XrJtr8dR+V18Mh3ufktnSUvcZFX4uNwGleapUti/KES+A6TK8H+oxrveRpcrE9XkYKJOoAHUOCI
iDvBt+RnphzpAr4pkjvZBRrLvDH7l7jnK/XpZJ0M5MrcsaiZpyWmRCzMoeKLk6v6x66jT32RzDHt
SCZ1hRjh2wskoV2GlR/xwooik8AruQsPF02ojDGsqIUPi1ZrT3ZjRN9Y1cwuj2cO2nyeLGYkLfKM
YTYxrp4IiSU5vA0ZfMjHOW5cJKoVI80aB69WCIgIySDf4mC6jbl9pNANCjSkCiB1KhtkMMcgMHZ+
eTBQZat2TU3Na87wNtk1b3fKezkkpHt1C2XJ40wX7Ag3+sXNZZipwRmBEMsqX3+m+bKyJ6eoFrs3
LOAEiAfwn4xu+zqo4hD/cvpvE7CN97FEOWGwl7IFcE4ja2En+BE9mUBGNe7VN9wWKX5C1Ji67xUo
hpj4+TxWw97RA7wRL7i+/tFw39HvX8KnbteqKaqSclDBIHugehembamqvWdTqJpqllt6TTtZelX8
vNNSrrabMU6ZNAB1KV1cLNsF6G0CSD5LllZpAFRJjwpeP0qKWRHi5zcInlUG2Rc2X68MnpoQlRFM
U2atYeDtaEK1uiBfR5+KONJxa0jCbkZW9WhuxpkD7Sruj+xZ9m/Bo61T4DSSsd+GGyd1aT1OoehC
nDn0a0TbAxsm9GvZahWGe6vTOli85cXQkhlIGZJJ0MytmdaNU6HTFjs775VcPK4uwJ/Ipzw40kON
Cnd0/cqoxxGyxj7PSv08KY9WSrCwDKR+FfmRd52I2W/osBh5/OI+8ebhCc2zfbPqxU1VXYoNLL0z
9FHCMfssnnWy80CUqV0j6lMLpFI+DcBqD6hXEkZD70CSCTA1a9dEEW10aTzjpccJTog0o23z4P7z
dIqHgemCLhMyKTfNTixWxGIopkcoYxDB7bF39riCnKkM8vp3H88NYCWxcaSahCjr4DMCq0b/Jo80
pcX6UgLMzXYaL/wZXPHsK4VWpJ+i/GRmq+JrGDNo4CwMyjBH2nN943hGeV172/yrbomCK43C5/6n
kVqJGDPA7dqHCuunmub15emdhAaRikcrewRGXsLO2FZdMOhptQABaC5BzVR9pWxc2SHUTS9rLmLn
iUU7yprmjl9EFcray8+G+hSEBkTnyQkNxTk5CRO0vKGUYfAKvGWGTigq7tpCP0pfPN+1ykIf+No4
6GrVg5fuC9FDhbXLnkx/TWJ8JjgSb8xg2Txu0YA5eRixdfno4o8e8mjKI+HBJUWdo6pBHkupamwt
RikwjVu6HdvxinOkvdn62HLDJZjwa1qF1BQmU1TzqQ//gIiZ4RStivayG55cPu/OwoysdiWDAanx
CNZwCg1008D4hstIwVgNXvp82+73EV/Wp3Zifu8NKsJT8olkpq57T9TDN/QBR+SweaRceW9B9gMD
uergXkhsR1JDgh+2KH7UHjr3qsCZayHNiBJX+qqWdb0tL+WwgwsApDaHhc2dfaCsVVUj+peom0/U
AaooBY9aaVw/6nq/2yqXRN2WBVltS2hMqCmEdHJiMxA4OPtioM5jPVOhtN0lGmDuOn8wJf+bY+eE
uHx4O9z9lem4MF2A5d4Dw9jQi0AWasvuMWwGJ6THGRG5IXd7GAn/TgyJOeLNIhnLLhRfgKMPZ7cI
0Yt0mCP3mL2atALQccQMsS0zGw5mntzIpbfsr0R5nksHA2vZwVKkRCF3kH4CwxZk6zPXURD+Q1HE
h+f90/K3ZMucwRxZVIQH77Gs9RIkGQD5OfqBfuodxE8j22V0GgV9mTQFUhnlL6MGl03iwhPp6wWN
AtTJeibCBx8d4khLy3SSdfej4HkGdY00Y/dDCbKqgToeJPKexprrlp/lPs1BzwFRpEIIAUvNjdE8
tpQL8ajbKeqMxwjikftFqlJLY6ofdnea1zxDCvADIxXjvAo3G6uJ2FsNg7XWntH6p+gpftrooqwv
IiQN8NAF+mXw48kdHjr1jd3D1MtEkVroBLE9fCPfHEPO57dyLm4uKJlhuG/eR1erY7oWUvRlo+2j
sd2dJr5UN1MSd5HiIU96xKwvi3QrMf7l2moWgBw912vJHi4IwzHP5I+1igCBwXZJW/OsTXs3OaBP
1VvkYrMGefkLkjs1RlC6/m/PAjFEplSHNQ4CKzd6ARvZvm7FaiHLiWR4xTi3Il7qQUPP1OMU2kOm
ydK+PiwMhJqr2+IBQD3qidW924/HRIJIKcW5JCkOzAw7v9qLWIh7n3d9AwAsYO2UiZHKjTwjRCFd
mSAfz70ecSbzQeUBjsePvlXxycSmXctA5lrGPQu1BARq+nZvFQAZPw7tm1RBUt1bAN1vLsHK06yq
WiKmKs9IJqM3j1n6kXbeZGQSzcsLuPurPp2uwzkVvQKxvdlkM1eQP+ZsXUyInSKVyyI9TK3P8oYW
UpEtoUGzzooCtfqF4OBGf3acHzt+L9OB1iG++KO1ekCofnzBnjc8UXvXv1couv7VGSs7XplTubya
1mJEniH/bu1wn7jls6oHrQ3q+zPDleTXq5djURpxG4960W+P3qaoWha2Ma6o7cOuFEP2SHzJbOKa
0qg2Gun4jkgqlhrQ8N2HhBx7WSUGqnbogENOnewZRdPxJrukXEizGT02e+Gw5/pEYvR0gVV7d46G
u70893FGamlLa/+AfcXeJKI3zmDg81XJmaVlsj+cA3jg6JKUrC8Kg7Z3uDN218bZ/kzjcDgBAAZC
8PED22nBQSSrcKG5lR0hNS88TW9EbgW06xDOpV1wsTV2QdsREkOrLhuy7hFaexlLmSNXgrrrLeCl
+0s9sM6i8A/AX0PrDdduotIezuLkHizOUPkBo8lIdiOD4XMt1OqcoolQHOGz1v76qVdloXnAn+se
MSMzTENMf7J64QZJdC5OEsXeX6h39mpH5JxI6UhICFT4RL/GC7c65bgVj1Y8SG+wXdMQWFRswFHo
QDO6Rmy7OYZTiNJLQJ6zodjopnakDF2x7tT9AKi/LD2/IsejFXBdXEuvlGrMpbdwIK/8KdwWHWfl
w9CXY8kOUz0Y0kuEEXxGadgwps2RcCSZnPCWYSlvpfN78ufOUe3f+OC7ac4LSHe+5G210Qh7DXus
OfDoFTctQFNlchElPkFfMTmJUl66n07y5zPutZuKRU8EpRFaXL0ZCP7V1gaHwAEZ/5uVlYMJyZ5w
s3WG95vYOzRr+ZD/kY7TicDJ1vaCtHAnhHTt73I0b4EXfPgVQEla5PxEup/9V6jEdYIxc44x/Kl3
abst80IiuPBKIvsgKsl0ff9xM0erooZFyXeZ/4EPJg2Whwwczduk1nLRWMCoo0pDuh4ZTAHVS+eE
4kzP8F4cHRooMKqlRQHMN0tRyw28c7ENDnyCJFjYXWxIKqKjeRKwOvTGmvAyuuFmd+6m6GrHxsvS
/spY2sKUbWeGyl/rGOHJE2D7gh+dcUiYmJ66gKhFgMn2M2WMei6ISCa/ILD7suAEHFuYGA6txzhf
TNWjkhDTXE2W1TVZG2ih3l5btHlepCtycMYOaVeUepZdWMjRQFxVmalbgeRFYepS6oYQdEPE7zWY
VK6Vh+nwgYN9M4atsej0VoLcEKmbDQ7JG1kn8BYr4EojISJzfo47yrU/5BxXjQYe3l2E8vj17lTs
ngs6qrFj+yar2szMojmiJjePfblBX1GGvd7pfNVoY8WmsrpH4tMaaYGrPSyp2NegNl7dGvLZqwDY
RoT3lj94lNNBqIwVUVPtFFFXb1xDB/nDHRFbg0sF0OgTpPOEOPOqOlnaKfZPiLnLXbLuJ6uB9gY8
mbujYlNLgR9Gg6bpA4qFuHPNm+KDyYYQtgmrx9H2kI5BD1h5Z47HEDeQUR4AGlmZd4sqMfreOUS3
e2bpGc31vDCY/J4Gq7i4V/L/PqNY7/aSK+S2M1GRNzzzpIqbFLuc0zy5zxJH1Aw+lA08/bWLi1T5
nZaLft6p2FJOBQI9IaJS1sUP+JOcJflfUPOu8Q4kiClmBfBL/QUC2ycL3J36XuLIBOTuuYgfBhbl
3QKJCFX9yAw0UccyezEB7XvMvSFDl1PU21JGEw6XN4UicgLJaX8z1pbmNjl6dYwzk2mGAa7CqeIL
YFa4WowvBs8HKk6zxy6aBh+HLWpP6PFZV7UKCyJWafVozq7otmvJw8y3Wu0ljxrdCBaqQXOF+vU7
SKBGDxMs4MrbyXOJAIVxYXBV7+AoijDYv9/yfDgsb9oZWiYrs60U0UcxIAtj43ne1dFUI4nas1VJ
NtNNUyHgzt07jINXBoE0HyHgHiJVYThQuzcmjfa7EMnPWsTw68J1MsJmVG+q6Y/BMjDin62XS6wJ
9VGM472KenImEUVbMnb5vEELizE0yM7xLHkQqKEX6fJvIXRszSyTnx6PcLBk3Uo9YCu1OJXPOUCD
htVvDnjCQ5kjOYeyq5CHBW+f2FsIklORtiGXo/zdpdz8pJx5sekF6HBoJH0Li7BnnNz5iQXut5JL
e/dwZaHU7lyahAgV3JbIoFwIPtPP3likSVkdGFaEXnRQFT16+3auRc9Artf7qB4o+gPpOJ96jdfw
/39r71CxTD+pATVn3+ZdATcCmRZcZISDnR/lZ6WIamQ/svbcayfPJZGuiwVcY4GG61k5iZzAdjic
LK+rXpJBFyFCj2v993JmJMY+iOkyW6YPVaZ9DPiJcjcDlqWxysbeoOngUwxeGW8qnEIeHzJEvcit
ugyM4n2lk7H6PAhb0EgeUx0XwjmRs+XDG0qIVrraAAX7cfgHLlSKqN/r7XcEtZeMMLc9qjxGXb2d
9mS14BjNzufq4UNhbH2bFGdERqHRH+FFlR4Sw6i54lpYfd/fjiyAvogVzrvGgfBCY9s+n23JO1c0
edmwjcZzTfJitBra4FB6mTHFthiVP6MNDPLAypPXE6W3285720gi5NbZlplLr3Y8Nfv7O+fwhc9j
Exjl4j1RwnPww2Kec7q5LQ8HW/j81/eMCqBwPRaY8BsyOgOtjfNIrYNiqWPiI4lJqGUga5/VwPMO
+jMFgq4D5zUYrf9l8hAar22zJY74/LnB5JxVw1rMghD3EGDWe45GeNAJJSbJ0KRkGTLYWJERPouE
sulasvT/eelRrQ1K9+cNyfZn4Tgtm7XUS07dszMEgWUQ2YUBoMVSjSqLaCrcHscDiA2EWBLlAcFM
/ZwNBNztwwn4L9z0ejxUgFR59AUIo2Bl4oPnMOUoj+7YsF3y3QKS0rzS0+SU/rT/ap/uJYlgqq6E
AyY3RYMYisc9MKrvUZzX4z9tVd+ts/5cSCYqpsyh4sGayUuUjaqCfCpCo04i/quCtQhVWDk1BWyF
RqjDvD47rsk1UqXUtCisnJuWlLWA36WTHfgZRhBIbyD/fHlkEcN0XABpeaUdlprLtM5vttZrTnEY
vt+mLZaxFZCNbdK7rdOYfguBMLnpWpTQJMBZQCt0fc0OTcqRGT88mHwND3mT4zqPVDL6kRmHR1jC
VhVZ3mF4gG53wsu//UXDu8ZFLuPhsYe1kKJhymneHKC87+vt3qu0s2++Z9zpKHRZcfBWB95/PVkv
aKdH6W4YRrxKHcAdJFhAtTKvFs0W5KIUixYbj8/t9cnnTP33jOub4oHyIGFQ5+VodL2F94EhF43i
Yk80XMZfFpeBYlzvrQ/PPlOJbT0MaeUKv3zb1EDUwt1oWhx7dZFfvP11V2mg2TAx7a2TLyLEx21F
lC8HFjgc4SwVYlmxWUimBXSHscaB+exmhjM+ko9Ti5HfGJ6nMXO6drVnxsG8pb0AvImFmkCfBOp/
iZWyNfnY13i9Wkqkrs/kODgfKSDOYTYeWzUVHCjQm9aPTfkcdmOJm0Usfu2J2olyhZytYVKIQ0ki
xulj77tsvI+kjMI60Kg77+K+AkTxPNtrjgo+DlJUhbq/DrMu+OqwQNlgl3rDTadue6UhQaSeRE9U
7zak9BC9j9txpM0f8g3ZXS9+Ln4PORjLbSKy49ujBbfruoxJXJu+VuDMkof9JjO59hrPc17Z2bSU
NVhritmReMaho6V3pnA/uUkqX4mRxE1a96fiJiz/EvGjdqCBZzrvXcaMKsVghxvVicUQDy19mFYx
2hzpuaPhxlccAZsPjnpdWbLUNGla+XO/+fQdrj7FOFGO0XZFXIATR6L7IkLnM/4CF61SzSw1odhO
yzqLHDVzbRF55zsog/ibaQfmuZY/Et2L5rorRw/wKF97aYH+1mXBfsCgzmSh5S2iCi5NnbTAHkye
fm4y8gNlg1/VwiTyt0NAc7F9r+d6PkbdgsA/i9Bb9plncPzYqd9va/33HS8ht2liWnWBfuAXRlXm
+pjtx8f5h6GROfAl/YXSk6cYT6Hh+ogGM1TyIoIByyKFL6uPxDocmj8L4DlEktVh2O8d9EIADmL3
+kiB0MdWLeduO7yftpVVhG0b5eJJ2iuAXN3UKiiAjyvXqraIBc8YejjaZ/d1by/2+nUqFbYLveYe
2TS/NBYgxdM6nW10urmlpfmQQnMQZhXajXCxHFhDBM71b35xZGjmxpGACY5ZDVSXuwUiUIvVO0fs
dAfiewPAK2pYYQhC+hFg8PXz750uBEd0nQxgeK/5eRRmvKXBVAuLVVQpyl1DZZpWeBbOHcM/ld99
Ur5jXjCEDaQJQlU0DmGhqLHN/V+Oc8OV0bYBtLr6MG8/b6X7toY2m1/2VUIH6gaMUYG4bso5ZpgE
hIbhxAwVPAAVTPVgow1H7pByMrhap1hdPxm1uu6hyJ3kf8oDvD2rOAeL9cW4r1HstEMX5uRvKBZe
XHNQ0vFOUyUGLOQT/6p6d+a5EbRhvwbWn8ivGpf1/ERjBJzQ2n7El2YVkfAfyXRFfw4NhQNJCBua
0C8breMwRzbGt1PrOEkpbdAnTGHM0/Gxve17uhZXjmIOjMPWxaMagubJMM8dOGE/C+heAHZDgxwg
ZPO6RSLbL8JiGrNdkQIqfo0e2BMoXVmUHDeEVIGD8euqEmF76ZJ2VhRad/rakFtBxQAWTEB1Iy5f
+N7IVFtDdr9OFGeT3InB2MVsGedlt02vRDH/yE4aC/2agBHvlwWjn7LtAWbcG3LvBe474l1EbYWf
PCsQiRdOX3VaXpMgiaqdM74OZnbnUfydw2V3DVOo0tef5dndbWfzRWdwv7LeGBP5ja38AA1uKV9A
qoAqhDuTtm4J2yiCG+EuwTwqaozsE2d8YQIykZD+PbIIL90kPtuGpf8/bszSHFSqCdkCs8yBOgUG
t689D1DIAUXuHWxuqbexr0lvO7VSpv33lX1i9OeiIE7U4LT8UKdUlTVMQrGlt069Xd7rLShcHdPc
dVt7N72Jg5Pbj56lAUIN2CtSSjptK+0Zru7Do0MLH1D5tCaKS+3SHMcqObUDEsKJ3oPo+DVO7agb
5TPjTtf2LCFvmQg5ZhKRHwGBnBRrNmJtlQGn9Tng5Jy8X2OL7mhKhwmp88MUNr0mWdkHkvqdR24u
AMR1U3oXUkRIyYiYoCXDihCEksO7WwCfI5PKttoZaUTMTskjncwG8h8HXpgTA/kzPw48vhkjXiN1
mAHSKRiLEvEB7ThC5j9z1LfdGmITyd1GD940Er8z1YLFEfaWlwwQ5imy5+sfQ1keQgt4/7TF/Fnl
xMAXCS5YAANGJJV2L0e32tvTE5U/ZbjGMrEwgOGrTVY1yXh32m9/RnUWvgsMHXe5z+sVzESnIGeV
o2P+sf1M+AfNBMqiMrhwJCX013MjVEC+ewKfQRJB3bB4qzcVr3cPQ9lo+7UESmRSifMss7mxEoz7
1DUOo90AhZndv7XbXVfdKFyE27FSlxodAworJfw5ukww/BNMiaqcmen7q4aTtr6FlxSZls4AIOHT
9xB4WVxKXi5yCjz3HnSx5L18J2TvgxadTM+7KOAdRwWIStQzJuLkzF6bhAaNGFTgTtQY+OECkIZW
CIohFkXKEwDJ0s0oyPgN5QMOlY1iLA2j5yvjENBzpF0A89kKRRYF+XmcsBOKeNtb3PO/w3n7hstO
m8ZVhIiQ9M29KGmvsZyt1+7JHFiHpp9Y2Az5CHT6wWepw2eTKRwWmrGmFCYGAF3xs66OGwHO4nIZ
x2ikAhvtqEB/Tfd08KTRqdTFo5LBC6eVSeIRghno5uF0xlmvfNx0bOUskIsntQA+Zo7ciNmTk0/l
Osj9PnXfqWWRdxs33cPxQ1BWdzfA31ipsbapHnL1ZWvXPiwpyjm63wKQZoJHyX2JU54ythkiDOL7
NvfRDzzEa5Mr+WjXsCpTiJKdsAdh2S08226XumkLBN23WqyHlCTu+iJCxUNMV8DYJczJOjsblWNn
W6MST4x8ta/DeSzCHVPxs3CY98gQyvmfnGINFfcCuL42FyihPqTA4+FrpOAd3JTc1acxKOOb1BPB
fTWSmv3G09e1FFkZVVmGNiSv+8M73W+rwT9CQlPcgCkDCrxzT8p7H22pNp6a5QitVAIjuHoDpywQ
jrO2aMRoPRdpDS9WlwpXMh8n0srGfElXffs8bQkQ6ZjVXxUxD6s5q0+7F5IB9nIVHpYBJS90RUWf
M8Zq2l+NS0ahP4GzrR93jMz/Erch+MIm0X16hi5/k1sK8/+/TjiBNmlR3NrUR4UXUvNO0e9N8rVG
qF4vUAva5jfwWQ42EtCtZkvkHEtkkz4Kr1Wlj5Ti+8pFAqyeYbnE7vswpQLvaiYQz6KWLMLbrhNY
JLgykOIWllYDhTNMIDLpA86+768TMComN4QHObAcZ2LeXqyZ91CCWXy5s5qbUnXVTO8FRLrglqzk
T7QUhpqk+ymVosxGgmFIoHn85KHfjrCRZfainaSPb9BZeIGQRnFZAdGngKGU+3zcRlTa73mnFyk6
0hqFb/vAxkSLM0GE/QdUMkWWsbUmbZNbnnlNeG1f/Bd0xgRGS0gRxL05XQJMc84uUrKNGDUvCTci
FjUIWzW7yDx59nvRHWK/RBPviZdJWyj2RBqHVVNHC9SpJNg7hk6tklLDsuZIpqY1uGhnVpOYA9A9
qUMiZIsyC4tF0uFQ6i7QnQLvEFgds27nADeKdeWxN3MpA8MKqm5ihxOQfzVMWTLCp8tTuvWZ5o/0
gxGUQIZ2TL32YRch7FCRS3H6vsXJ40duUvVHX+Dvz5ScwuLJk4MKpvjsTzlh9GK3B0dsO63aBgiv
2CKoIDg69Rf6vck8ZfkaQn5agWUBqn2GtlRXXzU3HRdEl1/Q46niY7MV3+6/HmVEco2qw34fKDc2
7+G079IHrhxt8UQ3g5IFnnNodytXS5XnKY6T2xQOx+sRnfavtZ9N1zOqtkYp0mjIOfL4CVcbZCnS
QM1GRnPHgUNW3VOQxVG/CKZYmNeQjrxAxVN8rJ3qCoE1R6b0NbD47FO8TCfk3UgNRjvrFN23n2V6
iF7xGfahFGMVMjshDlA2fG9F2VW948wPkqaqNeksVYfGSkhVRbKacXhL5mhebeRsRUTgiF0YRzwF
CZxbd+02tlr1OBJz7DM2g26N91l9AOtYfKtiCZFlw4obATLTcGlfhco1Yuai7JzrUnyKWXJy74Vl
i8meKzisZy6UDZgxIT3Pl+T4fvrk1w19AdfOwaJZxFq0NhvhQ+kdo107qocqa4WQwTlaHKdptypu
AltryPuuSRVOV80oUOnxj5lwQlqBquocEyXz2B9YpEv7vGRyITY40LZFokXIgm6h8qu4RpRpOnVg
5koKeZwaIOpgNyGRtKRyZcvoPXW/56Cxdq3Cfo7hr96ftclywLNkqNRIkSadbeBa+4RctpA7rFjd
lqscoYlv5WNyzqdUqKRoJ71t/4+2F9RnJC9Mh8okmBWrGixUf7VkmPFwsCtG+vlTq3MwL/d6NVA4
kiocoZ/+3gzIHfyBkP2n+lnGaSaCSKaqjUZHyE1WI/D+D2Tc2wPYX0D/uW/s9p3geOSUMcniH73A
EoMkJxOK8f2l7vNUYKiSlC44h1+fbLqwU1ubfUVWlsRGaxEquGvzQp0cdmwhRVlBKcVORgyr3Dkx
o2cUognXVkLZkBIyn8bz710Rr7o3k1P+Gx0DdQR4+Wi63aBEQYLADdJYPDgK0T4t9FLkG/5HaLcD
Ens1BO3uhTH+ce20x+a9GieXIHFfBvy62jVJtrUwcXjnom3517KklW0bEHBddrfg74XxWrmRyTOo
DaSP9s/xPlhTo1N25oTjAVElHVLKelNHfuijJW1fbyuM5Y0X/CDVxXAShC9atqfJBZytywaxD/rQ
p2lq7OvqgCxDIQMP9DA//fbc5ou03KHeSV+Wtvk3zruR7klzsirqmWtglnmAAv9wP3QibutWnpAr
KaYgj0PttPAlvPvzLHZjyuMJdtWs0Lw0CaXKXFJGe59K4BWXY5h/ODmWiPZpBm1Q33CFwXbSaSOS
XaMTA5zbw9u8MRTk9jzB63StcZ4e6O0gQ8szIZYH/KNFw3JACH+jZ3XkXuZgyGXYt9kT+Q37oMFy
0WzIh7nzi8IRko9KP75klqLTiFJBEKvXSTO51tdfZAZKB9nki1vjMyM/SaPsxX09xG9eNcjaBwuf
wEpLsooSWniFRdJRuJ35KiDOYWSPyZnkO5/k1M32KWwMXziCPr72PeLJdqDBEnvhcimPjhfW8XGS
15ZEzyMbN8RYbbMeeHIXM/2W05fSbSWYqncAbKs2Omx27ujDhnmevCrFGzTtD7GC0WxaU9eWE53h
rYgdy2htyl9uKVmO/b9zClv8alYEmmV3dUl2EnqxGNi9CdLhvQ8Q9Vsu9bZzqDnn1gtVV9c+48/g
IwDbNvEnjKRBJTVDnoGj2JZM1U6VrmDx8EazZL/9I4geEu7hRsYEGF72wYkdroeONORKjXmoew8K
EHFQge/gNzhu+isWyaIaGfJlttyosioTsDKOM+2JJL2nxl/X2ChXxWCi4gKO3Xx0ZmyVgSNzYnDa
bEVSXjoy/wzxrp/6Cex81VXfaB/naWHwHgFDP8I652gHBhZak2TAy2Vp2ABrs0smYm0Lmxg8lSvs
KNUN2rV3i+NZYrLrP78RNOpK3DhJFO0anQ0lsm+E+bwVff4rQmpmcl/dHK31+gnO3GNjOv/xcHhK
z2Nl1NB0NY5BElPYbmyLUh2J+Rlc2uB3cJhm2hyxmOXV0E3JBIPEvzYYzatRaF32FwUiGI93uvLP
xCjiZ82hbID8k0GfjBkQ5K97lmq3lXZMHRYKHmqyLgbK087BsMQ+94rsMGlm443nKuBhCxK9cEAT
qPIqCRcW1B5h76aKPAnozinY/S4M9nyQFhGXEh5SOBjP6Ln/nd4YnXGZqsxgt/jhiDCfJ4o2qRw9
q1Dw4eWdFxLMFtlbCaA3lN3s/L7KKLlmtt0prGH225EJGe753yBcXlKD9B4dGYZJvLpwpuPYPS/x
JvNFVniMOG/yf9NW6XpD8JeZVq5k3hwcHbwvu/jhaibPvppd9o7l6mFQt9I+K2j7RX2ifTvQgBbO
j28UKzdjacGusmDHiqQyfVbqYTvejpuc7+hzWvauCAaRvOpux0wLF6PVv5UfKgwZkSgCV3PYOwIL
aqwgluSRZwIMfm2qp3U4cvwp7qJ6GScY8pRgY1cXWIbL7fyPtIiKazrX/9dRNvGF3JH+XER3WPfH
+c3dLSQiIYfX9dyNVYo0B0c1sLC/qINHeQW56QxNVtwx259LwNDDGnK9QzegmC1cZlBFq4vIoRfn
6SEpY2Q21OCmcA45iJ1burH8Q684Awe0lGMXfNiz3Dt6LJF6zAB6BHn6fT1UhCf87nMZVo3/0wsB
Kds66LMq2EVS4g1Xw7SWnTOS9N/91lKvjrkc3HfcD2eLtGH1ZmBh1rgaEP8j7vQvu/IHIoQTLxKZ
7aTmQ2tTKMpj/th7f6DGKyrFu2jO46zbuOSmfr+K48tB5CelLN42Q0UAlmAcP+NyVgWC1E1ogDwV
UE0fXpahlhnH10rRVzzqgnEJE9NQ47XqiHwDuJRsdLL9TxIgj7GGtHYWEBOnYQB7JMBX/TkCE57h
AH8jns96UXF4dDXA/7jCqj28TAiFzy0PDMDs5A63QS5pxpeRC74wwi8mgDoczaX4huSjRAs8qq+v
OUvl/IWkqXnx3OcO4a0L7Yx2jKjf+oHa7GGFAV6tzfQmCVAzJNTYh9maHxULmsgB97KItEVcCDQP
3gz+blVsYMn8gGdXnuCD14cxxkjyhnv6GUmGPR4rJ58TXtIdW0bTLy9EMylLXcOeU4Crn3we9n7N
Zj2O8c5xP8cdZH6AO6ESgz9y8ZH1+a6LXbVXse5aBJGDB2gfdcSHb23257tJ/gePp87TrzgxbWsn
+rsetFpwxj6RoGUVd6QHb3ktvp7QTkh0Qej3zY4kGH3pgfGNvJfFKKipXoeJqmnYvGWhFlG/XUdS
QRR0E7ytlgd50AJMH+/Ee9bA1E56IRcMRFbM5K16zUS6S6A99aUKI+kG+1vg4g338ZL/i6vuVfoS
3YWYG3klcLoLIzfE+FmjVNqXM0G5in5Q17Ut8f+VpNS40I6dB7606WdIhGRMegLXiML6G6Y1rdpH
nMGNqqUwsFL55F+J+loanvfzNRNwhfDuJgDtpE6JTiHk4zmX5WgJYpPXHIkSXbOsVTpwU75A1vms
0c6/JMexv276W7hbjoCKr/DUEW4ZGpOwDlujoIW4sSda3TCF/bouTYC0qBhT0alNrEjVsu7N/gih
hfEtG5M1GktaW9OZMthX21tVl/vvnbCj86Tvqi2pVPGV+j/ZYaKhn7WtzT0qY1U4dMy/Loo4FCpG
vU490cVt6t6XXKgBiFVNNGc86lmy0vZoACtnr3CddYYOXaQ4R2T3i5rykQbsChETxzr2PNIq5OjF
t8QO9meJ39VGd6YAUsFWjXmZ7GItexnCRNHSmYNNifYYV2fcQFYr8KH9Oxk8H2pmevW9dJzrItwZ
3tmAlebn4+h+BzNDQyX3V9QjSr1+/X0cWpTTAIUoJnstRp9leaqeHl+ZhvJTuYyfyUIbv/qSAA7W
s7r7Wj8/JLYxu8iOiwu2/eyarCB84J+GFqYolMADa9Vc57J5sXVKycAGEZBBl2WJZ895urN2Km42
mjbTMRr4LEFzkdON3Jxj4bj81dcwJvlHgyc6hOzbCy9ftKjAjX5BOldiIs5MSl+vsErPpe/oQB1w
XtVdkyyKfif7wqD4Nq7ph+IjiD+gT4e9/q/PNboTKy/OG4DkQqeknC0nc0Fy0w+07KpVJqNO5yHl
jUBu1RYqflqtJp6ksSwmarWyUGyzLGEnUMI5TppxYfDyaIISKHYJoAaqqYhIimUawXD1bgfReyRW
Zl7yMHgrYs+/xbyMs6xggm06f+P1LlvbtF3JqcGYv6v+/BMYbANGqjUMhnEpc6en0Z8GE1SuFwe1
++/8A4d13UOREyMBbGu/IdvTKoxh4z8n0Wg0AUbK1Jx/dK7Uzh526qjDq1OyBlzoV3jWuZK0wSBl
3wEYwnFOYbzK1wtmpmQmdVVsNkR5YCcHqhqGVUOYTwSnCuBeL/3N65iGEXlv/nSmgA/yV3liLtM6
LJy5FQ+RlIWAPfVfazlpY/ZRGfCoRwPAkayKwwrRCuax2zNVDPDg/mGXnLldh/qpVB6JpkFk4rNQ
wj0b0Vu22JOx3Jr/PeQw4aqJWAtrutoFVLkRdDizFApauvKHVzlWHejhnfuZ4kNAH7UJ34axN6PL
wlvm3oJhT8LZjE5cyIcRqqjQ/qmYVFiGxaLxz6Th/XlNixbsYD7Wmv7UO/Y3s/ycevI2sPwyAWyE
pJsAZw2HW13vDg1Qt1FzOFq5FozK3Xy9zyzy4+2QoVmdaQRUp8VbyRJxnz4sArXRbGf1XTJHTjDv
TnEVSSOIU8UztD+DriSWZQc5f6fLhSMCfJJLtizTCSFnl9KYEofdsdVrBoef0wAjYpaPK+LlOJS1
mr59KqN83KLrlgSarfK1akA3LwaEJAUoLeUBFLtyIYRU5Cy2Re9O37/ZXd4EJR/g1tV22vyI4WYm
rtg7IWqEb9ps20uw3I/L/Epv7W+Uanx8MG+Ra/udpVYv4rGbe4MmKkQv4nfOuLlSMTe3Q4Y4Ev0o
yEaGUCD+0zY4euaPwJVyMAj2Ckoj9Zj067GcIBfJmsqFf5LRGVhUBV3kkeADQf7u0XlmxzgX1ARd
7+iau1QqLyNfaifaoOHWu2L4gJYlkEJoHe90LMzmV9+0rB7NTtkhD2D9WPMiEkK9HozrK1rM6PXr
I5TvAtOR8jDHQewCNgTet4pN3+wJPiWsSx2izYjnD9zwW8RDDpc/c2yZV+2AhIu6Dt8nXVAcH4j2
E7y0lL3YavZEo7lUdcMbwENBRAIIa8hCUAYm4FFpKjBPv7XCgVPTCCwOevHBmiW3LZzzrKaySfsi
+9hHrOecukXbEQFS1clLgcHDVDl71v+IZBD/sgjPK5ysjxyPxIhzTDU4ODmm2ExVOdosPJdXytbh
e1MSqLLtHVCw5wLpKoL1uusNBRc3K5Dp8X+ZRkiPlbE3gb0GeO+OBanYY0sWFzFwjFub2dcvXV9k
vq4KzRNMReT85TEFWcD6BRqPdGpaWtRUeMKV7Bo0d1Vd0Zrxzg2OFucP9eLkS0hViih7h357GYmX
1OGZ1eDNBShMrLYjlCuCRFAfjjTOzVmRVY6xg9qGjp3sI4jR5+3EQbDXT80TDIfX8v3F2yHZirFp
d/Q5VALWi/6tDpAvkHZG9bDQ1FTNZuyHkdXcWRLGI5aHED/X/tkIq8JDuQib8MbziKJpSvrFoAzl
coAXPrQkp3j8aMsHopnrGpEj57a95aMOe69pSXPo3EbCJCha3gDx7Sw/Bku9dXwT9RlFnhU7nFje
cQb3tN9aaSnw2+pfOLe1kIxOeHj11Y0fW/YDBo0JN+b991U/e+aPdTwLVOMH6GVbN64uGp/rO9Jx
EPsOA56Ml+CxQv/iyGEzc9zuy+a+wIW1CUJX9AZ2HiKHgX/Qy/+KhCXmkWNVV/6zwBneLNgQHmRM
aw1i7C31UpsbNOpcNqbpmnt42CqVaSaQFDOf+rgCpzscgMWdhz58xr7QvdNNOwGt9kDaGHUYU0og
uFZlvETY1SwRzAKkukfO3o3sMtvNS04jGbltjsq3uqDZQasHVvJsP3SHhXTgnnHPe3YkO4+ekxNQ
2OOJBbziF6yUqTQLBhBP2SIzzR+wu30hHrYv//uU/1tO6dBocXFnuRB4asmikXF/VRyyXK7jV6CZ
s5cIP34Vbt1He9ztIlHEbNHwrYXBkMkhvlBzfTbb8JqrJZlyLXvDv/hekq/fAnJzE+UgYcFuLoDc
o01KHLX/YTvV+OnWCmxdlhEs/A8G72zz8kaAdBiQxUfJ+gshxQgiiAS0MPtnJ79J7hK87o8p5pD/
8dVbQmEJRcZQ83bciMAFbEvI7ptxVo/gNarn7ihbttyzlKiv9775rKaUXjOrxK73K0JbD9hXLRd9
UD0fZ/HGYtJVyDvcSPyBwHsgqJPCAwzw5Rh3jQKoYRGRabirAqQb9NkTfDh86bN6zIRQn6giPn/D
T3zRzJMH3NVtdgbhQXskwxHCd2Gy0NkS2gIbwqGHg+YXI+p88Acu4bJhjgt+wrS44WZcZVvAqkvs
lht2Fw7Xk/yYKbSg15QeUY3zi6UntUTniP/3B4pdW6HIzrJ7j9Nc8FhmJntlGC+UKvDWjE+HF+pG
99VodKvOy6sqbrR74wL9GNK7oLdI9PN/nAEujmO0yTP4C1ProFaAU49xsZeVtwFzAQ77rCqorRsW
vqgyiwwJUxIioWuCeNk/yop3mE2+0MazPro09PGLUgW6XfmI/3tMF7eftKa3s6onBie9c+yycvyf
A+n+4KgNRXdAB8xdDwb7j0QC4QcjrEUl1mCMwInniML6n/JglU5HvHMUhdy0GskPVPYo0gd4Cir3
vLORqAcXuqTzavIWHiJRzs4qa26mJiQVqP5o5stKIP4GfAZyguJSa1AdS7DfGuHAg777q10zStaE
BCRSjbEFT18/UEEEt/6SpNvdc8FTcfPL9XLUurtLhGQSlhSm964vRetXPD5pPEV7quC1eBk2iU/B
EqgbwD3PSdl/L1PjvOUN6XwEeIRjd5q547g9tlpHdshDOvSAU8kMXTiFBEaRpgLl9sooX+sltYUQ
Hm5jVkzbMP1sUpr95B5P/6czpiRAEv88FiKU3GKviFWFgciVENGwPaHLoLOHHl2TdMdQUbL1nMMj
G9fi6x74OOITwv1+VOhcfCPcTwvPVVXgjA+MVXn09ZVqDCxnSc7aCvPMCT8ORyR1ULR3XjB16rTm
oGiKh8b3t4gtmjKiVxHfedM0O0KEL4xSLf3PsN2MzRc3Xw+PzAd1ACRCcHKimMeWXj70jCxB/SKX
Q2GrkyqXBr6u4Q3f1pG9JWvwELWo4ALIffI8FKgudGbIc2jLh1KbqhoI1jCamSOSIyBfRe1Unnyj
1XC5ZJ2IyiyCkQyT+C1KmUiU+s6lhkNl3t8drwD0NzMGXEX11HOGxceHqTVuuoV4cRt+ujgkceiW
tkar+SeaiHV4ApVXoebE8opDsBWjtcRPmvPqQSozXVh1xR9xJdCgM3ICzl6JG9rfXYQ8WegxUY42
Qz4tKgVSA2gqvqvF6IlUGiUb/E5fKNp6S3Cn4fDaeByfvc//sgmbTPsWZZ99AK+R/ozsLtWXnHHY
ChIV4wgfIcN5Cdz41eKgmljBuDouSrjUd6oAvQND4/X2ynrCYUKJBESKNxuqLTpzPrv2XuBTjy6H
TgJTBbuO+4H5vOXC7Ra6ZzzNPzDNu9MGsvFHWfwSrPf5ZDjLNPbIaE1+ZsJCcfEL4kqDXo7aXr9Y
ERyLYksZMjAJy1ljYl/Fl0O2xFvzqLi7lBtv9rG7QLGYCAKt+PVvxa/flkUoV4lIFpRTyCd5IZfb
2PBBSM0v9g5vi3NUiG/cSO6pxLmKI2M0mIidVais9wdtzLCO14EdJfrUf3A+Q4PXL4AR/6+R4LTe
H1sI+VH3hhj606Z/1/f4td1ikW4PwvrDsiT2z3Crh15goNL85uKG+WRFGLZ0erQIoZwsJlu+hBi2
GZnFPwGHK/pfgG/kyGbE+MyaovIQFq9RT75GdiYrqC/K0qORvd42D76Z1I/B7Kh837V4nQr13aGZ
daetZ46KOXhSafsPrnjVVz7ezSyvW6fQqkLPBtxOlEm9QTa42f9AKkvxNJTts1Ku34nDNwhloyLa
fhf4EFdNVxQfPi/+blS1qjZcB0WtVA4kLtWV+HHtab+I8q8GtVnerJYezQqRTXpEjs65LYLCMa1d
wuHb7Jjj7InlPKX2UfUZOBdJZW73L/7h4z7iFgyWxxDlZb1aMqo/ybvDqmvsuk9mwm17gM5P7zzO
VfwPYjivTB1df9+Bs/phvVgTU6W9hbtiy/+xuaE0J+HcdeCk1x5s1qRF8hdAQib4SflhXFazSMPK
htEqC0RiiQcFkL7QG/ACca90e185kNlDI3v13xnIRTAkDaF0Bdu1DZILKqKc3++i2STDuC6IyzI8
MFZ2b/hA54IncjrVR8RohPPTDDlv6iTU+cE95RF8XaO6gWNJC9RnbaSokTd+IRhMMa0sEYwXKARk
6ZBWyF8lH3TyMOg0xmTx/zrDcJwyJitskNWmmA2Be3J4WyfKkCMCiR/kSAtxXZZ6szXhGhdL6UiE
nEBu+yZRostK63PkMj4KZHYOhhS/STWib0BOfjbU32I/m7PnAeKpaqln/p7B++b2KmAnbQHxUyf9
mj4Yx6AjgXuYs1Q/MzRnvoX/QHB3Isvd7XHhtnckDLp1V+OvzQlE/kr17ar6j/GZEw/NJF2yyeCT
6F0KiTEccjOR+F0+tMtM9TQJdq6jI9AJTGOOzS458iHPgmxbO8BBrOvi15/br9GQQahAI1thpGRP
0DCVsI4snaOgt54J0bOAvAc3z5NU4hUFsy5KcALBm9Zmt4aliJ5p/oPC2L3x3xk26GnM4BX0ECDH
gg7CmgEw6eQskgzEX/TlGYBcZTrPwxbEFR855rd+/vGrm6O4yktUCJsdovjtQmPmFt0m+ZNM8NQ9
ksVmXmXvkWiVqXMcCiZhKehY7+ix7mZijaYTm1TmE4CsGfuS3meQMHgLZlxLmUEuww80LeUH5+Ge
el6wUY53b1p+baECHRtI297EV123qkrn4nsAYaKG6eloAF8t4HULk1I+0VEBwyvs9W6ihN4c/MW0
wolqWRrQb1NQ+uzjVU1CknhDZK6Zt7dnmys0C41j8OaqUamFNkB1di7dLftLHORbnHLgv+8xZ4YS
4cuTGVz7Mr+D4E9HuoHSQCBI6mK81BakG1eAbj8xjdi54ow/O0Kn+rBhZJlZgOqpRjxVoaGpRLP3
Q5laF8+FRwI52yAZLuW2Xi8WSIPrp/dsYQdJHfI/moT8qrbBfcz3Xys3xK7ezzpFLP3Au10GOiLL
yCB28eBNGVy6O+FWy9ZiOqRczYRL1mz4yYF7zLzX3aZDF/707eWbggi4ZjuPXSJtFbBy/DblI2da
rbOb8Hgm7W58OeKdJ6GAQDNYDQ229+/LtswvtvQ5pQOAWQ1QXhnxLlDqwmqqGB1VA0KzBi0RK8YB
ENs5ESUc+XPG+91GM7pYAoUfCS53UheOSLWfpvqJhqaCv2OP6lz/g5pwDTFEgiE+SH8g7gKrMHmX
huz9bnHv8LKMhl3LPn4LyAUNDnpLgCWf6cVjGfNyIvyqcug6PiAFpA03xNv2V00PrWJvkVckBgwd
Y9DGIR5cvGlU8sWWufGF7mbcXIx/zBPtgj+O/8aP7CrsJQJ0u3KcxKrElAXQDh58gGtCMAokrAMo
5bCcvVTBOQDmif8Knl1Ncspl1NbLKC8rASDuIF8ZDn+GMASx1NRqlyVYi+1Ma2AvQmxVKKmGw+x+
78OEyGIXVy/p3v4KXPicKMC3h0GbvaKHYjEtW3fBV0+4frG0KcMOUUXiA1lwGULK44Rk0I3WMpa0
obWZo0JlppoyFFHLXyH2VhN8/U7aDpJXrI0T+p7g34/5Lc7iY9poB8GYwzly/+loVLExg+1mw3lQ
70qywJKJQbQYs1PgoyBTb3lHlz0ze2WplxhR48o7uFbkn+6JSos7oYPnLCijwOaYCsGRCAytW46P
1UkuOzudgD5MUTSbZZtHXkwZ6nCLALXy895GbLZ3jdEFNX2v3SgM796VqfEYpFrRUus4xSrbdknI
hB8zYl/YMr1Q727PuVgN4uZRHnXxirFN9j2wLGbYboDG/ebASMFGexCB1U5JCk2b4Zs89/+djYrB
gumom0v7rGdllS/hfBEmkBGFG0D7ZIg3iRL5XJA2xN99YIC4O2YNuvfx1kLvYMCq7s2A4vqUl6KE
Lp72NZl5cpVbR4RedQziJoM7lzJChZ5c1PTUnHOFcP3y8f+3K4VFFnD9A0iVnGVq3UY38OV81qSL
3Q66wftWU8T1mAU/ClkAgfNP6F4jPRtpQ3yBHTYzRXmUwPdBOo1v2/1Cy1yvn2IFcFjhebN32RhT
hK0/wf1pGwa+JqZIn4WhNNum1pxutixtBKum+yYD0/y+qdoMNG3jWvLwB1G/LPhoKoCypNsqE65E
dnin364sPoqZrFNz0Tz2/5IupolzHZS3OjP/8fVoMEzhcJUHgmuaASzaTBdfw83BdYC1zFOifVgY
DJx1CpGWJ36bG4oBmFbUgMOIjUAcCltwp2OithMlplwlWcyYBPfppES+m+zupJaKtoA65uOWR6s9
yZIhs5Nti5IK0X9k2Jh7VtWnaFAxsFOT25RXB2sK9nSb0osd1aqxiJqnZtNWTiLj81nO5u52iLlt
FHroNL005bHeKvUIFJHvJmjKNNaB6lCmPyPfhSFKCcF0e3xdpvL9oNYd0CYpRXyuJnErMwVt7A3q
DyyuRT61Fw3r07ZS68kCBfdFUyQgoHAhZfsmUc8/oIb/887pqNTBguaaTaBBtpEyqdV+AMdTE++G
i7ztCRvBy4kTBCNgjaAn3QDc9GHJOzAaOgw5nAKZZdMxrtMaT/Lw2LOg8DYh3wsgvzjCCRH3dKWz
msythWL4KLk9Vq9lUo37AC9BypdBJxg9DUlescBJUbe5uwOfudGrAce/ViZJFoDcB7/NfU7WDfEm
AYTLetOYOWXxROeiQKS90KeySIA/icYwX67fHrr05edwgnYAbW9eOvxCBhE/jpZIkhfdpDuuNWAR
UwzpQ/7vJEVJ2XTu+Z3t4f6LWJ0tglKwqPJpJPELka9+y0Lgx8TPQjzPfJqOeuJDfa9/avl37jQ8
GWErx30TvEuLKb8GEBw1V74SzB+Z5DGPU0oOLLIIDHD5lH3rgsF0S0GWNXAmkLCBAUacoA6muT+6
BFzneFsCtzy2YKtbdRmom6hzqz0riJjbXvUcRo3hynAn3/SIgtaPOjXISz9y4MHLR1WLGZm7bQVv
8UDeTSY/u7wowcL4kQbTjknzOzRqYQnig9c6KfTw9FwmEsUoTXJP58j5WwFUIHY1kswydaPlGhH2
RY3r6AFQJJL7fQ1YUWNItBsaTJN5IB+4PnRQTs6gNb/C+indXZTMBSd5mqdBzvbA6pP5upUCnusm
2SXkLZ/XZZIW3QLcjTnY0aXesCmGlM+OJxHQqGP0GoAArplt8a7JrqxW6AzDYJ6SHlz9WVE+ar8J
FEXqH6eBGh3pOsEn3sOXPJ4MIyqYtbGf2OmiUf9SnXpMS5WQ4YPd4h64WBGU/kJdV3jZ36dH38wD
M0M7HkKN9JV34+zBdFj6GkYhEyH0HpKFXMEVdMQcwUcWDiRdleIrDy5MjljuQSCuxkV6JKhP64dl
yxbNJMI7S0VeskNkGvPpnQYWSGXf7SDqG2amfYhmrjeLCmRVhft1DOytXKAvKwAYJ9m6AAXhNwBy
glG1XYfSozXdTKpVe0D9rTuDREfCxEi+f97NBTQHbGYEQdbGU8BKi1ycaJfjUjoATk3L9N2mJQPX
Js2I9bdoeO7kRhYrPOU3TPsoZ3s+y2phOGonKVtkBIJ/ZojAuZkYeE1t05RbH3xZvf6K/Y2T8yUV
nD+OR4RUVy94VxHMxZvmDyO2dXlxuKlGA8VdUX/wvaWJCG1BtW8+HMNFuXtt9kYBf+zLgixoMyK4
UyfR9fMII5UHnwklORt8TAa+HfjdBJAqZ2zbs1Pw91qczd0nhGORVtDantKqqGw4p2o9gPCONrO5
CIrUW7CyEOKMxo3M05zLZ51mRuLYGXqXK9FHvTJjEwAH82T6ZGHVl5yi7m5W3AQck+gHF+wJGkFc
rIrogmmClsBgPBCAjYm0MySBHQssg5dplvyR4rmAXwThuEMeHVjIuQm2nIQZXcBBlH1JdhUIeQA6
LB+9ePr6ihN1YjpDb27raYHsQIajvu6T4+DkrZGRLImPoOovk5b3J1bxcngDKeRwp2N2msF1Bufc
7wHOzFV7c+aof+3iZVS7yzUsrz/FLvuh+ZFYzLocElixt7eZes4Ywl6s6BeOOxb/MCgsJ3uzOP9N
lLwreOviFW+LLm4c9i4oiAqEDcmP53/QgeM/6ON99PBzZTJMvuvuqgsGDeky4bEZ5vK36AJExYV6
PCOKcdIEcDrWgVDNxGin8Q4gdEOLqOjHWwP2ZVW1Jvl1YIsELHlpdplMUzESEFVvyVNo5TkKAahX
F+C9Wv9Z0vDxwuk+uITE6+muM4D4tBw9/Kz/QU1LIQyVrZZpgeFKYpBIT2ln51avXRgyFW+SbSD4
SlfQHwwIRLrel6uROnk8ayUMqdK6nX+JitdhgrwyxJ5M9GN05JkhbFUD3JWuw0omVxPxTrtmnvAk
0SaquvIWrzCDsu6PFr3McoeiJWFSQATKDE4ShRBArJHYda9U2gAkpLAPzXzS1XtoR4YG3TRLlWLm
y+6tuHhIOMEGsw2qGpTxXT0lKKfUsbH3TpNsJqkJR/jQ55dk+ZXbAhw1KFXIJgjjNc0DBXjO18pV
8xGoVWpJV3YeWu2iBqzGMnYiwXnTKpdhtxioAl2744DxDmnuII0fQtZ+hiNe3irxkM1bcRO+DKqb
1B35vOVjRpc9+7RZE3JnG0Js7pv81Gs3mgDxHcDPjEqxa+mPXsEPILn9gO+Y8OuZd4JdpLqHnKgs
y8ENqIyXuIXQQagB6maKNPxx22ujUORZd/JW5PSJ91RTfbIjbkgGiGes2gyjpVO7Y59rcvos4/cZ
tdlefzbaCt5zLHVrXODpi/PzJkY3JdIHQgDxR5+oy2rsXIv5CZTnE/qXtGQZA/uZ89WIvi/JbRgg
3EAL1WSIOobjpUwNlhJqlTeA/FhE7CDSTCJaos5DbT8NTJRm9/EGU6ZQ7RLhBYz0sbx0hcjnXz+C
X/KFEo84lPFoYaE3nJ4DSxlg9cEp6NYio8PPlmnEn5rZZgdbLbgLQQlr9bGczLtu9l2EOv1Tpv8N
q4j6DrS4vOXoT4VTLT/SsQhsaoasYBblday8SbCWBWcbPENWLpDOlxt1sXSAJ4buUPVXm2tBtSDD
KaqxhUp/Q2GMLoBQfqDL6tWU/jkdwOydACiP0Zj51RfYXbu0aMxMvAwDGmJjpzlqPDXyOAc9G7oo
5uYqZEBMzZis+Zwsu28toDTgV3nN7OIS9qxonGa3d7P56oFx/RU4OLp3gXXoeXRXgCs0De3gADpG
xyAuxBMtSxHInAaSlanr72bBX8VY//I8PkedeIeDic/Ek4ULqo/8D++G2MR5Hx/tcvqgLsd4qdVC
hQVZGZvquiNz00yxt/pts5q6SoYDdG9eUeQiScMe553rTdmnh3Yp+YA6/UvC61JiwjSKAjIg6PDs
TzyjRxa69tiNMm4EcVcyf+l/RXgD+A08NKXrKOKWLBaZOG6Tie0FBnwChQkMfdj8YEPnmzJN01l1
Twq8uUJy94YcuNmNQZ1VtzGzsxCDCSq7VMjZJ04/D6xcygocOBYNO/JihSjwG2XWopy6hb/zj+Wv
eu0zmuhd7aU4xgrXgGrlpdBUUWKHrbyw/Q5XH065dFRAWqQUHtlIbWM78XXd+bRGLYWAAwyNia9n
4Qcpr2tuWfFdUaS+A4qWuR9UEF3cF3VYEm3wm4hlhNb+7hV6+rVvhXTltk9ci1SuG81R1bnJ0qU8
p5jQW4AYcP4UcRSDaoETnMJ9916uLWEifamQqFauu3UxRVYd7Yh2m4Y/qSItrZp16CqY7U/sr2gQ
QRHJajEoCyxJlE3yVgbl4jIM6IV7dA/imZOPa1+1UHwU+BICbTxBtpax+Z0TpzymUM1N8JDEajV5
9OfmwHwzEx3EqlJgJj1n7Qa+V8F7r6jYMouCzsVaDp2b97JSn1gawBwS296eTXjoQvqRz+ayUxxw
SKDmE3KkJNY3eda2Y0S13ugGZ613xUUatQqEXb20XzB3LEyC6/8WdOd5BW87Sw/1A9e2w1mpshlO
zR3a92vGo3fI0meEEretj+MTVcBRhzzxGBrH0iB9gbkBINqdNcSdujBeuu8K+6nMmpImo1Fy6l4L
XusuXaApE64sXSq4qk8DDlD32UGzfBAF1qXR4kpCYXJd3IRpg6MgByAq3Kt6qkaaH5yljQcJWcXo
qmb4CuZdhgFPdvU99PfIsT9/F04vkqWXrKPyceeQcnAykXGVIp/vdRGQS+gaTI/qdnrhOUzs0Chk
N6LM5Gi1pEAMxatjTN2OviL8DGc52RSgSU68uW2I3NouNpk/ip55xPignF+9wA+1oczzf+U5rM3m
pzDXT2MkD8lvhUsY/Vs1VkvMr0hpzgS9pgBqp/Mqq+ww5hT0NvPfvNF83MgLS7+fnTxejen+2Xm3
v97gdIh7hTdcvKz1KyGCtHtlUdiYzBfdlXRDFH4Pc1Dtk8QDqR75moRpUU+H+DHpNlNoD0OHq6kV
tCyIFse3p11BmX6/EcuRVYfnDOEiPzmHBplDtE2NRlFGLYxp4qU+ZkVYK7uNcHpMVGmE0A0Ojz2j
R3ceRgfWSp0ZdZg67bQvvtL6luL7xsYsQhZUnajJZXBshk6RF9C8lgXw59GU+3r3qWXkEkT/Oql2
nG518V7HJkyZBMnbZyk2mHPzvAFl190lGpeVlI4OauO3wI0CFBifZolEtuViPEzVdDN+zLkxy7Q0
gd3+rlEz0XRK5PGLWLrsqhU09hg+VAwJizUjFce3rlGPWr3Liyvx6SmeO/9fBLbbTaVkt31GYaXu
Ez6PJprDeBz/Lywh4umjnsQ1UccKbEmwyivC25uNJbgOo3RI3OHFxXnmrUc97YqD+k9fvneAAqzR
l34xwMsmiCFKh1qd+AK0FDMrqkqIbcgA4Iegwpdujy1Qx+26DDzMEpgx4ZWZ/jwn8CETjjkJsXX0
henIx3t+9msVkWCl/pBWQazCYeF5IC67aE1XRhjHDYLUq7jMON1cOg/2IYwLAWbaXovCXpf3cWNF
Dq7F1XEwNP94Gm9CxfWr/RnT6EnJMl1ClW3/56EnClO+VrT4TPSVtAI/22EwoQOh4Eew7f4aF1nP
A/CwhTsczmIQMUs9o8H7Xd8Mkp9k5XPQlcL/CD5SLU/cJ+d2jfFHtiJvQ70W8MI10gyTXUJRXpXe
VYyzix/OkdocWsQ8SkgH2EODDT3MUIJxM5lV6X5URX/nZmq+kdHdm6dV4Aa1nqs3Vtv28K2uV/uJ
7GE+Gw1DphjjqDecrwpAZvOE66PdDeKyRy0XAYFAJtDA7UrXSzFBNkMn3G9RKD187/L4C8ucY1jZ
54w8/soUc0hICQeTxfnGwzXSMgUMKdyBzuHADRngoYzpgD90SFdxu8ozmg90/118xPiYqi45Fpmp
YsRQOfCEpNH9Pxbb0JfyMjmjcF4fbfqEUgSee94YRmzvf44NkQgza7GH+vbvTwkG5iI6IG4CAfic
Qjw2SPAwbz3m9hn6DySZ9unXL9NX7PAu8jTMbzHGvn9L8sUhj96KJnfjXMIjN1mBP/GTpEnB/1D4
1rJZgoa87QwQWQC3bPR5BxE2glbb2STgBHy4PM/rNpmH40SY5hWxsvwI7U/kBsVeZZAnrcilGfxI
nMsSmbshRrbWexH7W799IkMD9e5g/mMf1xz//80sGHlr7Y9NXWeYJ137rNvf4ab2eeGcB94S+DrL
zNHRKlRKkjQC+iJNlmWMe877DI/sTP34eKPbFRHw60b1YaT/MdcfQyphlwcbucWSb6nVaUSkD2ek
iWGftoSYlu+vjKOyWMquWbzTbnCmmmZE4HnCubKhS1SDPFLdO8fRhH4UME0mQdbw0MAb69n+2qYn
JV+rfyExoQiUvVyQuHxh6gSi+uY/PxFT9ueY8ODt/JXtp2ApyQ1isR1AK42SMRmtz23VIonRtZCe
IeMBWEu1f4/bps1dsCAF2PloXMAyXdKR/2FLjAo3jvXD1AU33dxe0glFEx7u0Fu3m7kWSrRwCZGO
DYFibVIsI+mikIxIieAZv52N/7bmV7Ng6w7kN6cQns1lBL/iUAXInhlrocjd4d9oO9/GcZuaT8rk
otc2lyPHxyEY1J/iFpi51LZWcqGNabpGSMrEFzQSKyPABGjma+iJpr8gQya3PwNPov59InnHftWF
8xNjZtO4OlxVhi+szw+Yy1LEEyp+Q0HValRI8251nv+ttGb/IH76lw5M5VlrGvm34y21/rEQscy3
NZbGXgqoZpci6DvG4r1aQfn9+uOrvECubpee42sX19L6pFe/jKsyDk5W9ewFNBgLByUBwLERSKm+
KfBRPgF6xI4cx1FvF9Fqm7Le2zT3C8rFuGLHKU3tEhpAmPatKvMFP+GxHU75aW51FwgXKT/uypfL
W+rjP3Q1qamqJlMjh4BlO2cLhVLhsQ0WkdgYgd4eJySJEOXFIMCIouArIbQTih43bIzVNeRYFJwN
SbkqRVrfyw3rem9/Tk0pzJNHLg9TsaIBgD/pyOUD7D/fbxSQIcQyYyfySSGhj8lSnrMJTq18Yd7g
mF265J1OiS9KBX+pa6tosGGiORgBBXklt6DvO4ECScWMi4PzkmfDB/QDPsR/rQN9PNOSbKuqMwpg
aPNyRT9FUVlGsKlYBo+z1+yWQC2d08lqiDAZUuOr2CTJ3fipixAvDmM9wP9Gt3NrI5QaMnz93KUj
Q8WX99Vf7UIt0fMCvZwDiorYg5AucaS9G+iWJGPJWTw0kx2aCWjzibjgY1YP5ooZPVJ0uBdi5wkw
jBGkZ2fHvLMyazgNmOiy7GbL5ybaBYLucFdxgxqaToA283iYNWsKgfADMFVlMx/rHAXiyI+Cgzkd
8cPcm3mRwRgqRMrVLTZbmtSVIe3lYEJ/K2+FlD4TB/Qzf6hbOksPvrnHvsBax5/uzC7B9KEjWFoH
CTnonVVIiGIe9G4C87ukGtQfHw0m3NRzrA5rvM/0XcVm6zixIiVrmQSU1xQ/ds0cMCdYRu1vBO9H
H/Rb5XH0Rmp+5UwbH/9NpDt1EKH74Z0y3g2OhdiM2J3o8kvwSc8re8AmMMVEZlOZ2jrE1vf+O/hz
n6kNPn1DaT0XgPu18q5FzYjGuBzoydNn1wNveMSS860E+vBAr0DNz9vFg0wkEKrgCtHqfC7kIIKJ
4wvJZ7vVUyNK/JA4KY+iwwty86LmYkY7iJ4vU9OdWxCFZG/Zrt0OOuvpPrCO9dQG9ObJyrlsaxgB
eJo1sgO3043CL57iUgDgQwXL5kG2xN1zZhHy35enw3euA1aGXXWcTaVzns1tDE+wX4G4OI/Trn4Z
brqqORn+2oJmpCPBzaNIkHqjLviu37caiMJ0ZwIreQtxhBsVZA847nVU5EyTNgRcMv3T/upquB5D
dOfRZVsv8qhXqJ7Gj+AQnG3jBUjXPDKNeSaU6hkCPEYc3L2AKJgJC1RgO9ClOWuiswnbPfepHwOF
cVEidcIjLPhggo84jRJcOTU0r+qRq0bTxCm3QK6uMfR8zCLQcx8RgYa1/VJcgJIVzxwQWYc3kTSA
h1SmCxEQHomfKlR97Jrzt9e3J3v2LhMEK1Dg8o3UG8LugpN5iVl0OrnK9De8wlDXer0Ck6ec1kx1
jZm0js69tU06x2TitXo+DjdT2eGx0t3Z8arfKhf5gyqrXG1KwW7NBJtXwglFtm+hN5RkneYA2NIi
stf1AZM2EsoqzNlaGNzJz2MHoB8AH0+NTwtrTIlPG1I2O+GL7aVdHewwmkt9vgk49DGbhjB4PvBs
pRIXXl87To1nMsK6dlpyo3jEmLeDPxz046vSWT2/KReZPfMvTzT8BDxvCLdUj3kr+6Hr+SbZI1Dp
NrdXxAw6su0ZdKy1D/SKEshq9sQFP9vmJjgnFqmYZviHC1iA05NsTlqV6HuEyuodZzmbx/FNbZMU
xSZBwj7YgxdFHTk2f3X7Tq/sGusk5a5TEcvHn4wjqMszpnXE21dcZzEXx66SPwZJDti6n7INUuOL
JLaMQs088tNdi9npfHB+ojXb0KXRZKYkC3OxguS2twyUe1a4Ltq+bHiKc8oKvrCvsQYliy5pFi/q
XT/B9A4nMNXoU8QuriufjrTjLP9HFqiUH4vjC3Po8+Rtbd1FHqEvBgVsyEoo0It/vvPa0LTWxMly
g3iB4cUNgmxT4bc7EBziiBeWKmCWz41+7q/5PZHaYNOC93oQV3GyD3AJAVB2XhGwDTOoThfDQv1z
WtwQXeJkWeRU1Qd3AzmTaiHBDsOyYkHtKmrp4cFJmEyressvQfHzQORU1Fz17PoTBHdXvV9lmcFu
AvPUSov3oEl7LgC2TKpANUf0c1I348g4Yckv9NZTL5xYexQmRulAx/GExRMHMXYrR8UmdT3Iw9u0
2zMlkNtMaJp9zjBuxvXbIFf5ZRfoZ75oOg4SoYs4AlOfIu3ch7AHPZRBgb6d5cJney7iR5XCHyji
PiHjEpFRcAbE8zBQvSQkwgtHivsVYEBP/MVtQ6pnarYQaysFLr3grRYqs6+NRfL8tLQkvqAAupPl
r3y/Wn7hIuj5U8Q3E11iscXX+aGIToClts4T/+JjVQKESbA6kq5t+s4BVJprn8lAUkn2L9WcJSHa
aULTQ94KldgEdS4MXziDKz5eusAhpIaqa1DwjGFBZ4sC7nP+89PrhGrkq+cLAafj5G7CAEgGqYDr
MzpYKvmKmNJnnfxbaSkBKu1AHEfS7Mm6MKRKyjMBJA3FghBij6jQHz8HkFaoqKBY6CMaRNPMKvIh
/aiDxPK2qX2BuFzOyD/2wQaNp1P9BKfWN2xD/CUSLBIBUW+zp73NZBoLCkMkY47CRJB25t+Cjd6n
p5bdY4eNTGINwSrfWhldSug7QPuCH40ofcQRvtiO38HUPGhx5uVSCS6Tk7grCcWllWwIOuf1hmva
UilkudE26nyCVbGemZDCzHl9nH9Hw08yfalQzHd8qQ3Zq053v3aCDL8gBsmSqxOb6whQxScnneje
3vEor5L84nVTR3/IW0AwQQMo++1LhsCECo75BOde04YiHah5CApCJCUazHT6UbJgIsypk8TQTZrU
T6kvPAy3keEsWFqJiow1S3y14IVoQ3mlFJ+YLb5wRCxEgJNCT+Cb7LYxLSNA+XwQmj0ktAj5Z6TP
7CEuQQstVT3i4h3Iq/xTS/f5Cv6RxD6K7bbzkiAc9X5yRClb2AJmYzC/eeGWDvQw/d7iMTK5jIpj
6WUaIwqs6MPYO8yWLfPH4Prmoi32CsVwv+68bfx7iZQdmNC9fpNdI2XZydOedqCZkCD+PqwNEugh
vkdKknre/0bDWhwL5EEE6ltfpI8OE3ToOZjFwpU1SDmKT4qDFcGl+jnoLgeIQBV+c3JtHvIMPcVM
UT5ssqMYxuNAQmo5fuBaXPBfBAbtlovplitUYH4gTwSUGSlNL+XF2sL0Hf+R/xO/6/DJfIkktgE1
37Sx3DQSMSg8Rx+W1aMY+gLR9LmhKY3XWE40fEPXsKg1ojZI8nOaXLuLzheIH2AkttzRk+ymzuiJ
f/jwqL4vKjTyQyHhmVlw6ZnCUQP1R5sHiLhDHQ1hkjf7gEyGiPBoPOH5vYeFp7w7wyZPr78Cdzzq
6b68ZO2d8/YBUDEQ+QELrlJZXUZJtzOh3j4OmWEhiVNLkfxwjA7h5uriZC7z4bpx6/Vo2pnvCLNi
hokUVAjQtb+UOBwY5olYX7V1yxEfy6W9NfRv61G6JiRsQtroM1QjYutWMWAG6SsqTtamynOHSCop
MA98Csi1swee/N5TpdCSBYFb3hniei070/6153yGpUP0AkUDecaBi68SBMKMqf2zuh2Mc1LwOKTm
mNDJW/PYOAHpvuf4MUJcXlCmimPMjIDZRFzws+E2Fi+vhAWfZVydxe8wRunHacfq5Lmjsdduvtte
zHaktW4GQEz/nogQLO/Aqg1IJbXVvCwIPyatFnKkyUA6BE0CUMMihHTo5x6P9KQ60TAPnkfeYivU
lxKMyFvKKFBZuGomSPZ3trQpGl0lzjSFh+Kjy9Ht7Q+nIzbxwkkjX55MXnFAOi/8zPdAItFZJXlZ
8X9iqpUIMBbGmsHUEQlm6Gri63AVRRvnaqTGJOP4619Nq5YBZ1xEWn+k+eizeLizrE8Hx4icNtIt
8HzWD/yzbOcwdyyPIgIy2sdAK+7rwuwg7lXugeQ6d0VWovr1pi655nh2ZnK3TAyuT/9H/2nLVmBV
SpBRUGLE4uECRyPEck9d3jhg/3+8jLKhsrsy1JrBzynnFAgJrqEPtSecnQfXPDY5AGhPIFJqeMlP
/EZ4m3wCScyal5r2jxrVmzjoWAAxvGf0RaTXm5ihLii2Bds1YcjJ85KfNHVDaT7kB7yHe46WBG/g
3igWgcJU/QVv2C7MthHU1JJN4LTQN46U1RaDRXSPk4o6DxDNyW5QZE2GTjeVNbADUcey07Od5JFW
PB+/oJ4ueOkX+BsvhG4BcidK+c9o03gk33sNNokZE4FGZ9Qq8IK+gVSUf0EzBYLxeXISs9xbc/vV
z8Ryo0wNnhdPHZbi2EeF1gi9mnyb+GKcOaAEfp3+bsIsPxonj0lp+eE18Fd+j9UjPfPC3VZ/Jv1v
XNiqEBrXrElrZbG1glJL6DaChXsBkJ0xQXtR4Htl0bvXTog+j9GcLqSsaUEHE56mjmxoMFImQOA4
WYRwbOsMHQKdURGBS6lbMNDxfA1eGEEYdI5bKBpDMzML2FQlyG7jCW8o2wJ9JXbUv+YFyF/0vNAN
eBv5BgPta4QcmRsqeqnXcb6cojhxdy36T/loj+5xYyZOx59QY/i+2QmpEVmYIZZC7stBQVEfAUiF
hs4yFznkgPZxiFmWxoDkuTjcd/iWc3PuNdDW0/ek7y4hm0ZnAp4g+v43aiqaYoISXDsIis9Q12uK
S2fhshimFCg/fY1XZYUn6ZMWiI56Nq2UjQLUn0B5dmPYYX3ANJ61vZXf7RJzST4PbojFgW2KYbRX
4H8MIShAxH19lk/BnmlRADQHw6PMHYbSXl8/RnFgoSqA6TOijOcZ8N85zqDp6Kn+Pnzsl/Kdxc79
SU2RSgE29elZS2NStXaPS4lzCRtPGoTcSpfaO9ZQ2AP3R33TFRtvBA6gs4ml0WGGeTnP/UIBV7TH
8t/wbVmLwzvIJuYYr0dqgXY1/DYXNnuzm5g2TkHMnc2N2On42azJrr1QzasOge9S9zWtUwvVE/in
OsnMEF+NqjaQk1s1fEOfpMb3wwycSSwFySQXQ9pVARUpjB2XguAgf4e1RAIxaLrIJvfVGsCFDXys
KpLe3w3D68jv9s8BzHAK6IAwU0IpZXOaDjYn0OMZGoyjkLH+k2Yfxa1OBrMY4K0TY8ezO1OdSns4
Vjn58y6EaPkuf3H0xgJS6mC+H3Jr8+bFJEF+E0dW6UfjmZQaqadvZxZXhkw8y6OzN0ZGeYi3xmEm
96aocCWc4cuOzXIdcsiGKx4UtrMKjUZUxpzBf3ByhGeC9MG57ZTaAK0raGvRHFY8SLUd+akAEeOF
QLoRKexNrZwYVVEyAj+rN5vytRsk2FtWNI+ykPoNu4lwpp9Zo4eAn5t7eZZSGpIyGbfO7HUfUpcK
SSF8adApFwFR9FuGMjCTpib6lVJEy0Ip4DdSXdobrxyZG3M/aTy4X4gFrUvuf3K4PuNtJ4MZcHdW
Ic4V3zuQ448TD12yZqdFkX0SUSi6bTPZlW0jM+dfPpYmfgagNzVj3sA4R92AMAXIN8K0IlewHDdq
xbZVJKWqRJzXZPRy50uy15mmFuTKy1LkVLj3nmkUp9dDzA/LQw3KRcETDA8PZvTWzL+c2GLeEYZL
Cggo2k5ID2upEQdxzgmFwTcpBMW9wQ6i5XlO15SfDOP2wh0jwONzUJOe8XSh5W1yhEQwrsgCjxaB
GMuK4pgf9pCtMDyEhn5rak7F8JKGQeWCH9VwvyH271iHq1Q01IJ8pWGkSI3dY49IpBUn0qHHX2xR
IXUr0vQ5b89Wyx1xOmDmtXjkkV4zQNkNhHXzqXKItLoc2T3c8KN8rkLbockG9tzuPuFbZMcj9aOZ
qJ2/fZQayESX9UQ8jS92PkvJdNIOuiKGgE138JIVnRZdAWlh0i44V/9RybBwIMsCk2rBjIjKLnT4
279EUKAjPCnRQLkMlrr7kca6gAisOFKLvDtDuNJfnfHFvBhS1+ivbhcVoHNJeV6AOoPM18qXYeqj
gg/PaDNwfWUW+dNxGl41RTCYb0U4602z85OYZsZIfFr515+/sNHXiWdVKHNAf2cFhakm0n5hvNT2
u3iTJBZNyZFt8xaSwjOv5oQ5Rt4Uz1YrDyJO1nEvZuXejFn9MQwfj3cHdB8TikyWGzsb4yrOnTia
axbyo8phAt4PdJ2pDriQL15HmiwJIwDInjZSAuCF7mBlpgq73fDu+mSlxQTmPCYmgCL7zy82Jfrj
lWjoMuh6uIEffEYz07rZhuksnd05YA9eAvxVx3sms/aLmNorSBwAtpx8aqM5YEaIbYll+GAVkPaz
UQj1y1vTVh4d6VYDD4Ldz4yW2wCbBB8jNO5U3jyOw1CqprXBfG8Rn1z5EnyhRUu6mE93/Yj9KmVR
14VYaHAHefmBZvQ2z8thZX8uSaQs04bWGk+eMAjMoNDaB+4ts20VZh8j6q5RVzu5wXrZFKni3djg
XWtfEcdwi2V0ENKKeasT3WvW9t4xtgTrOFf0AnIPDcycNeXFMigcwwNO8xgi16Xbjw0ZT3PXMM16
5pYeOOL+x758/DL1b8HKjEIBXxvl02BgDstvZ0F2GZEkfDHixln6N112+maxGEbmsdPu0vClhZ9l
ilLm0h0wclVbssZaMwMrlWiu0wLci+8KFfwDt4GKZITegqyVYa48IJrDPqH8iyUuFNAurEzrI2BP
RxthC9rTwzI7S6tOoCFDsn4j7cvHHwjidANjh84VBs3cK/LJcmrLNSNqn2GMA3jUoLu+hU6zMnyq
U37KLwuU6JB11N7df+H3+bUiQ38GqgMYOlXopK2eYdAlAJXhO93RLju4l1CMiO7qcRyksbhnFH/+
nXtr3MbbliL7ENQYLSgRavlxTGw41C4hI56qYIY9wDvqNlZ6ViPoI3pMTyfZnOhILBxIBrHb6hRE
kuJMzbLYpzWZ+/WUZPpw1vwtUiQjIVGVUkni1BBMbNlekdIi63sztTY/TMHqwgoH8Xj20vW2ZNK3
8DPvMF9kojzKEXySPOkCOfXVAzpu34FFEw1Mspbeay9Eh0QJhP8lwI6ykVLbSqTzL9lZsnn6LTtU
3XsPAT3bMxcRpXxQvvN7Q2cWlBpe/rfZ5wg9UpuHwp2+LP1B71pLM7IjfERacdLqYRN0t2HcZHaM
5xwVEno5XERl9zWGT+pmtObulFZCDDVg4beSmsYF7VJ5MJHMXk8JCO40LCqhU8j4OQ0xU1e7S5At
o/ga13/UmEJzXcbK5+PISeYFIsNTMZ5/9myuqQ4iiY+KiA/WOWBXRUnHudvo/NcmVamp3JOSWVVS
mkqLvGiq5CRSolnnYRE4hnddXglRlaGj0dh6gggjO4cDg6snQhX8c1GVo39IiQzrERqzbxlSComj
xfJUweyjwwePkYQOlNsSVC96pCQGThtd8fzLihf3YTb0vzOIt7ed3b1uH/vAN+i5yq4OfjpjQhmz
i1MYpAdYK/vqsS0p8TFywwGwMEIAP9EuZKr67ZvlUOUCQe6JYqGsGaQCTFUAfzx1/IGKgRXwO7rW
CCHCZYrev9d3bHhxsGpKQ27O0kKGLkyw5ysdMazAhT4TQ2Chdlnga6NSvPHbR2ArExUbqzVol/yU
oX/VNLSVRkZCCvjTz2KSWPAISTPplC6aqY0EA6fVxINo75Rt40I9jc2gphgbIYuUKbAL4x6Us0uR
XDOFru78hrCnW1AaDhwXQILk7ePjj85Tfduzne4xHtI09Qj9YkbdWZWeRW0BJ9xrY6GRo/lzhqE+
dBW0Fmm6MZzhrBP22TBQWLxxEZxpip6QZNr2aQIxVoePyYAhZJpoy/fwn+9rbvcxcFTJsHMt84+X
CtC65z2kvoGVJ1zBI3eiDnGmvkuc1/iUjgM+8MJBkHhr/62pWZLqCb/DE5eZNSa8u72QeqxWfqvr
UUTZJQhZV3hFOBGrkMb05jl3mtgEV1OuZTtqFupO4T4+hOlxDWtxHlxjH7DhUSwwDq7etrQ4wtEA
Dl1zrW9HFd2vbIhk6hQvbMbNF7nYCYpcY9Dt/KeslzO0c6Lvl0W7MZbr/vXcrQOZTOdrOLtTea3a
a2D81B2fDbd8XI85zFaH0uLFYfN0osjDYq3KPHdn8j26seKKs43KVP7Plotf7RJUA1tQ5JI3RzCM
iyUQ2uSqNYMgGJ96uSYPIcFTaaC9vgEE0efJvcl2YPVfUpj85JdoPX/aZ0CcWrD+YR1FX0wjQJJa
rCTb4jIdts6YnWV+YkkRvEiZMr2duFN7IMKHwbDqOv1/QP7Gn3AfDu1HA8+MZyIRDvKAw2/TuWF+
71+b/tQVR8iIV1JiLHwsgSUhVqV7AbxDhx2/WPc/Hg1stca3Mfia4I5sUBFaTdz3Jj37fC8nPjwJ
47+Wm5Z/U8DpBp+57X1Qq8uZB3qObAps8hWkni1eh8Ng9sODtanxMuqVnLS3+65p5NDjmqc5wKWz
JoHcW8t1Vj0trPi5yzVVT0AedBuZhhv8mgZuW6/7d+saAy1g0//rzwgq/GbRGwho5cgLuShIP3Iy
iydthbAXwyrHIO3caFzdwOJ92VVFCEm4rAR4qvhYNWS2eWokrf2kHsydb6nTjZXBcRYvlEnBqYC0
z/vROP2P9/YHaMifNPbc3Jh6Lyqvf9jt1fFQKS+Di8bX/vXGIJ4p2umthUdRhVYSvmt4gzofePHi
WFwL0TAH+aFwAXz6DDcsfTeepLdx+jUD968nOyMr0jW/f4S5G2YuZqCvbwBArR1gifpMUAF9CkYt
RQTNy+3Ex+GjU8DU2TK0+TwFzpsCx1ECxYvjtGfIus5rYqjqT5qC7a21Vqd/3mEROvG1u9sweXdA
rSPIQyNctVqsQXsU5eZweZKeeHF77nfjBELnoJ5LIouZ65nubtqYpGvONOGHiYzkQzMZz6BsoTOL
Obp27LmM7OzTyUOSBn1ZB9Vq8yzMMa687CGkOmtqf685hgg6s8hujK+q45vdNGvTfNrHtBo3a+KZ
oVofAZLEUrOYr6uATzYk+Jq3H1ijntLPnvSzwP2e9uivr6pq3K9grHBql+OOzwI0a6FIL22G8vR/
tUI3Ex/EmNhmbFdTZecl8y74VjyaV8oRxjA0h5d0pZcM0u6n+SjqvXb0+T+11xJSJVdRRRai0YiN
fv1c59q/QKgwG+ja+/UB1d/Jurvc6B9q/heImHcRJPYpZk2tdwvvk7Xd2b+KspQTuOHReVabMkEY
jbroq5LgOZtk7v0V1UFX2R55YCAG/i8wQhvPnZ4nrD9wuMLtHosvVCNFX9McF/GdUnd73S5U5HAT
70Ic9rxlm+Q/dhS9EoDlAhEtO/GNMnkB8P6ezHYVI4UkVab6mYvMNcMowLxaROrTen4nPFKnD2+r
paToKWnBoOOAJbxGSbA+1DTR5MY9AsMDw7xvxJYSCnRulq6zL1w3He3KAgeoHB2h6LHLUPnc0ZP4
ZTntvIgaXAKe+SYuYbGEy3nfB0SKJY0MErNLfE1S7VRZ2XUqm8/nCiuR/9KSE8dW7i/O/QBAfGKW
Ucua3NuL2vD5HMhA6dSL7ni4EktJ+nnOubgHcPyYvhOXvyf3TEbD2yKFWDf2m4QYAN/afiucxnfE
oW+QfLYtFMgoFuMY0J5OnIfzZzzKDV2OImyULQlCGokMnxkdYbCb/gJeyrqdZQjAP4RzCLtHv9FE
3agAR7nTYpZS80WmqP4krzP9/zy+/E6cPqYYnrzE+S1FjI9kgue4tS2OrR5uxHmfKoEVGtMMqWFq
V1mPedrb/cQj54n6KneM9zuB1iFkY7TNcV+PrNhEz8Wu25F5mo4l1L8CGpB7niuNiuZWTWcuHFpN
mvLOHVlL58UBzvvesqkAqVe34/tnQ5M884MhgM3IrE/SxBXOXorz14gUArVdKYHLlxtALnszbnxP
ErJbBej5V+K8vHaBk+/D6G/3PeE2j44smxnNTlY56jyAnW0MJ93tbl/QTSjEhQv8w0WUZiWlCtAw
MJM3uiGliYJ2LqlkO56k+QRN3xCNFLPifF81O+ZQKv3GMhtA3Zn8YCrgk1fcizmzhz7O4WzE4FK7
WFT3CIocTu1lIIKfQyDmlO+RN1fft8bFyGdcGWIuNMzZdAIVJs5Wd4ITlj2MEd7nHNpc2yIJtQCF
eZDcNohkWaBdy9nCXzWE/n6cecsb9BOQWvjPQLvbAhpKaZoORJ0+V9EdGorAXQyqJcFpWMUUwqjl
VdO6QhGUHg5It2eUeGF4jyC8U9vq7cDx8H9Ozcg2XGyQrWachwpYmIbECy76M7SVUJfZqVQ2CQXj
F1v8FBfH5K6rGHxYd/kioQAO1GP+qmQmVTq0KSkNoTn4/1LLc4RtE8euYkFdj5z0jY1pzETI0TuX
5xwWPoOl94X9Zc1EVBCLPkEI+8JPOrD+h735aeDDamgwbB2tWiQ2QWAenAcM+zCgrPV5a4NKiYet
iRF4m87mHdSFcXUM0CqbxTEqgEFab2kE+MprXfKu7CSGikl2a1sAvKt6S4aaERquk0zvx8CQYYDd
eAKACd+Y/h70CymlYZ6dfmUq1UG4I41spqTIoaOSniKxD9MCQYXT/RPLA/q+ZjZiCypgrcNm1bWQ
SMcKh/80lTVfTM2SfPwedqulsEBFCSGCxk60l/n1D3xUhrzEvhgmbjZn4fZ2wxQ0/Xc6QV3irBD7
kX0jKhIuKzasCnrpQmJJ3i+GjMhY8OkwTnWIGBmALq88UaACl3MuRRPRLNYP3EsbthfHcAl+o3Gh
R00EuwM/6DpOsUrb20QvlqJyKdnvA69MsZdpaxRTqq1odw9VxkoPHOt+tRFpBIdsUODdOigWzvS/
JvE71lao3TW/fP4OmIe3Vg4tIdAoI4uTmHG+UVO+JEp3VdmQloyM+dIFQ2/VfaTf9xVKcNWyq1hb
NxykBl7FEQQ5F4oBQuDq/dOPbmcBJJLTfSzQOs05Dj9HOj7/GU5A7zmT24+URZWJ2hxyvuTaCjPB
IS1VWZ0vTX6GjP05krvilzwvD0iWrl/jgC1dprFT+bCP5/rDHRseYu5x3ElUNRHkoD1ShaKcFu0V
SalN9kd+1jr9c11HjmmAWiF6scqle0GX8vhja0WeZGz/18LhDZ3oZV0BIjGZIUPAXokCw23lMN4a
HY+haJiAvWQLfJA+lDkElCr71lqRL2Rhu777aDXLBEgdSExGQYyDd9C3zrlqoMbfWUZ9wOX0ZnB8
8RdISE7Lwy8ObBTSKMvXK758FCTPXqcCbMBfOjJG7Hdu78VtygoQNDCyxwB/6Okmc91igofgvgKa
5ECpIUS8H7kFJkoDbXu1GyxN+rySKXtyBkPBCF2OBHOam8nV6Fyp6dl/tO/YLfvKkKKkO5h+6Xsu
ecuBEltwjoCrYHNNaSKSVURmX9KWK9cqMOOu3NACmOO6Qr6cfDA27hBsHPeEaaBTBSuFBkFpFJww
5exIrAaQMNXkr25GpGX62uGpxBN7tshvv+MgyQZLA4hEJow6RyNFDOMOei6gXsgfDoCkPFzUniY6
OwzAWwffxq6KG8J9zoOXxyJ40l398vWrwihZtZhkQIeY6FVBxm1OlN9AKOravhsYlAzebXzu0/Gc
51PiaO9oSZ279plsqiuSPlMEExLEdYJW53o4z0C6WdJ3n0iovWwkDGKAsY5PJyfC9Q/jTjN1u0Cy
2ZR1x+1Ww2pNyjm8OePJWq9Tftnid4KcxoON97Xq/bh4zl+hk4fa3XHanDqsBKI8swT+QEbPOrnK
vq8mEpx9zdX5Hm1+/J9VKxuSyvBZNZ/cBYYdmOh5qGopfsNMBTb05IhLjwLKhWJn5Z2bmLBG2h8H
KCoZVxGdFpmGv1xXzm4ENTh7uvKScprMEMOyF8io4axtvcWM40a2FbfpXrbZ/k7FrhgaS0OxdKlk
3J6nYeSu9D35cnhUZr8NhFUHgISsCD2ua2vet+xT52Lyxt9szrg2nf8MSQGx26CfX6YrkzObx78Q
59UIrbfGSsF1mB5ipeXG88PwtGnuiW34k5Y2SG1//Mvosgnjkxk9Tc1hhYjWYkgpztiqzpEkesO8
wJhd5C2IIxVcbVlC200e46wa3onB1pzG0XXjCKZK0F65ivP6ZbyuuwWuFCcfqHSFx2d06ZhAib9u
EJPeSB1v/ogxDNQVrfi/YEYkE2wt4xq8m4ey6v5ukDvAewnylpkEba5OvGcxN8dY0q7+ujDu3wVc
zM6h759tWKOof2OvdH2NxzDg0O8shsOMaVscpxaOHHZ8m2y6HgFTrQLQ4XGjlqm5yScXKLYuu661
JvvsLBo4gM3pkaMH6ItNYw72gnJg+VsHfPv7Eqd7OvrBD5kfsJBKd0dTLWRjq/Z6PdepszJHCFac
xfVvpQveI4t00q2gM1+aSIiqNXVKq7GRDiMvFKv9MZrjGcGxBsLtuTASj+IzGXhBGKwogKt79mAR
FbiWm6AU3aIAvzOb3uAfKvAOkVgTOPgScsVPFzMYaZupvVIrVlVVc3FahAZsMAFPmmkib+uZFTlG
kP1e7W2QVSJaUZRh7xf2Aai32T6TZlpavHSGCELikSZ0WaywSt0rOTWpPu5L35UHHOcp6K7uoPz0
+qWwSeH1cUnsWkjHmUqpkkNQuwgOa9XtRvGX8cqog6aL8/zFmWXJK/VKjMupSAVELnXnc2X1v9IF
hrAchpifFLZD9VCkJBT9fPcIuqTgpFpLmx0Oc6iTUeH1LPhlt8TFcpR0j6IrtHBKS/FzRiACSPAN
KLDOuU42ROByD2UQI831b85nuecGmbTnlmQQ0nLjZYI/jdomeI8TCTmVVLwncARdcgXC+PUbRaQs
0xg/GkCK+VsKV+w/i4HZI1CW3Zno+yTeclRVeHmVzXA3KE60L3tyOrvz4YB4OP7oAYFqTEnakZP5
xslOcwCcSRFeNlxDNUlYhku7x2vJKVTYvD/q7NTu41ZdxASdpOIDce+yyMRbIWT8Ktg7kGwkKmtM
maAKjoICp4lMKISZJ0j5vu0TSp8RCu7zRb/bUvkBqomFJDy8Dkr7ljvD6uMRD8mzfsSQtYGWzn8t
+Vzi0eAbL49CGtmkbF69Je8M/QWNOnRtUDltNA11a5bn9d6LKdPLNWrYEP1hdlW0TKLQbG97gDk4
KczUCJiueJDDecF2zZQyhEspkiPKwuI6hSVTUhN10Knuv4ldBZncuiFEW/vNKtKNAkjPIG5LUyFj
c3o9G6GzHYgKrV278yBOeT13Oy22IXvKp1syP7VAdCfIUp35+4OG5qrnnDcoFHT+GUIyidjaUKJH
6gaq2jKwt7RAwnSN/mxJR4C+rrxinFDNpQHmCG3M7IOKqQY5oasGz0rl20vGiz8XMmec7MJg52RO
znvqtumnPvQfSSkebB8y3ccavVYoTRkF05Wz5T6jSeZdBMVvTNpykLrc3QDuEX/c+J+3wfkSl+HC
MI8iayJ5hUrWIKmjrwZC55hrZmcuNN5BwY+AMdoICAj4L02/+Xy8fHp+C3NxeAbBwEZboG0x0stT
wTVeTrWIp3fQ/e3yG9GwC4BtS2W1BU2NCW0Ia+P4S67KYaqWakyoIKb8loid9qs7QVtGjtEtPWZq
IYnR6WIr+vb0rwheFcfppkUoJfpJMbguY4DAcPH+RKRuDu/j1SfIoou15z/RC7D85lNoIXEmmr/2
74Uy0ksf7DdiPbDw9V1yA6KOuyMqKTYQalj+M6rSza9c055JOJo+xRLJGsFNob076zEAComShxih
pt9YH/1KwEit5Ac+2U17rh6R2BTgvsfcAf8Hl9bog2MHt65wpndWpQq4DlF0LhZKspsVo9uttWOb
p0deYtrQxOszCfZwaLmvwTCxeRqK+tlepTa+k7ljQ3s+tMHYlkwjZPBfozIL5VxCqx38opGpmtmu
qfYCTgVqvl6239vgdXG/eYGocBc1J03bOGAJzfsIwbWYDJOavW/I5frpn2AZK+WcQ3fqRC2xQCPb
/1YSdU+seGRMGMKBN7t2gMuw5S32ICYP5DirCQGu1Ar5osqh4ggTSD66DNQ8kJEDb4m5mldGCNNq
a8+G9lBCOVVjQoH7e39DWm3I/1Nv85fwkajt3h59jQ38wrycJSgvZXYFgO8YSvNu+MbON4yqwhWL
RnV+d67Zcwlpte0Z9QPuRHS1LDPAa4qPE+8jSlGmrVTF3H0igbBOq1NFRtzGza7Q651S2LfXLYoq
Rg7kHyp4IWWfLpJ65q0Zp0WnAi76XUQ6pihLPOmO3RIqGTHzQxWkw6MrH+IcqBto8U10+Xtf1Ir8
XReM5MihW4TQSCRV8HlSIAejsna1Snaq1zWlMUXvmtl2WtmmTwWG6pYGaf7DXKGN8Q7AAFWOcWji
YtCgyRKEtbVoUI8SM3VNsn0BVST9/5t1idqPFozG7vZixzJ4aj4cJzk1zI3Ei6CLm56U4ES6XjXh
jmNCZOPx9gx7l5f8x+DPzHGYpE7q3DtwyvMJmcI4rrYP0KgE+KWSwh5RexgSpabRXu3AvXCJ5IjH
TfPQ3moovytCfNt6taNovRHoy3zWra8SzsQL115PFmzKpu7qx9sOYhcA9itzflFc37Jcn83pW60V
cBmOf++bu0FqJBJFBt4LxP5xoAn709VciCuq/EaVb12FIOWSA/uX3qpqErL5wUuu4iP1PxyUOPOH
awES79ezLBnY2OkxfI9gay0kxvib4A85DGEgIXNOTaS1RtYDhs65R2l37nzVIF06vhFwm9SjVtTo
Ljbua/Bnl/TxHNk400MPCGlI12NTs1av/bvqFmh/ujl0sexWVtrj1bU+4Bn+jREsnzq9zGx5QuF9
jyCCfrw4Mgg8znSwdfphhOLV8/uuRTDJN/c37w4tddArayDOtaRWMbGviGJuarTFUTx1ByrtUUzg
fwKJMHr6zLIaFcPFZxcv3zxIH610S+WQDT3f5nZwVzuZVakPMyiVzE0hJNUSi2itoJVB8w3RVxhO
xhZjhFRhS44W6h2Cbaf5iH+9z77k1DOkovwLBfY7NIxPVxfL4F/t/48EB9RMxbgTUDrXLPUGEQyE
u3biTk2ikvM72WCzCH+GKd29tGEoc7diNqHLFW9FNHRzajdSWRVgCIWZleNrbiz9XA0Xs1L4sAZ8
DNK+9/dnsWUcF9y2O85CC+e71KzLTgUM8Lwccy63ZYsoZUoAK9t2HIfOkmvuxsyPiwXvuRddR0iR
3HZM29iw3wmJy9eWWMuOmEhqj6qSAc2F0D+Ji9gVekDregnHlgMBAR56awnGDfmW6ALfuKo/El2d
yd3d0thzo2hpIu3AudP48wNILBpiDdkreFPTb06j0xHwisLyDzIfbE4n8/MzMYcG9EWW6xjT7tB6
HyJWAbQt4rU+cpfcP+a6eJ6XDK3IP1ysA5sadvfPsHXAt9uAayVclANtLA7ki/wbcwIMMhdFxDVo
upae9d91fHTUwVxEiAvQtvz+tPUvuFUVg5f898VftMHwhmCJWfginQsxFGXTSl+GzdFIOMGckixC
jZ2nIpz/IAnzlz5xVLxJx2+v3EJHG4bWLi6hetQ+vOw3V2lYjD4pRV+kJz9MLmURrFY/fuuduLgA
VkgyI8t22RN5xaO5jlBsHXLBBhMRl6NxjdFFud5blmdAONdrPUVIU/XaO1xhfJ+eplV+Q9V4d4JL
HbVcfCVOFAe36WODAF00bV3525VuCZtfH32oztnPj32gkhzu51QanXonGIHiTjrnJoFcmxM27hO6
wNa5qBjBQCwUDlE724HRxo4B0YM5xHRPX+/Sr0TnMMwee8HMiaBP/cLKvo8/anx8yqrQsuAXj60+
TlGSn0WzRq7NvF/989ELM2UcgVDPUTV02ovTHpUzWzrlzAO8afOQL+ANwGQuiWPIyuiRncV0uspW
Dw7kOHI25NQcvPRWOsnESmcaaSV+ERhixZximkHa+Q/6fjleYSaMuPPwXAik6xJtdl35eLqpCbbl
H53tRH/UfmJ8eo6mxpsoC1Ty36pSYEd6N2xF6f2FjKepAtqIc+18AlS4XfQs5WgYmQhMwmL1L2Go
wLt4FQTj/E9TQOtu7Xg8HYCqRvwz8OsxWHbzmKMSNXprI0Vugo9Wp/mKLqAXsjBIbjSqha8nx4qO
PPkYeEULcSUfK/q8UFfYV0KT2WX1aHb6IqhPDCuhVMCAeyky2FGVE6s4n/ipfXMkLRPT0KXdtqG/
SkK+yy4M5RUN/RcEILiT+++AgPFN+8QRCi4KyW+SXEHOUxoj2NymTOXYjd1Ec3arsgZoZ3SYCap9
JRP+qvLwTHz7/pSHkQQOCb8q9ySbpJCB8fY3Ew7zUwZ9nrQwGTizg0D79RIdpwf847QED2YAApn8
MLoZUUmUPIgOe9mp7u51oMjTwXiS2KSEK2QFdaBvUvWSRfH6y2T6tbdvQ0eEsAMxgOdaTVPT1Gwq
pFwCQ7EByy7UG++oUfSVKYlCex7g0k+BqnD8WqfdJLtvAx3jPD05l864rvOz72HnB3kbKI2O5qSA
pOLJtzvx17GSbFU6BHMoHKKeydz+8J11GuObxfhTIxbhdOgm+aIlh0PaOvWYZZWAAIu4x6AiYc11
pUJCQGEES47vwc/1OrY1Ndt8ksjf8qx/eYJSQbbGLCePBLrsHGEMq8hprGEaAXQf1NWJ06IpQPc0
P7WQ3zi4Im/fB2lDk6l560OpyFHtHKDWygUjFL2UmVbvtyFZ0knZ5OHDzDhH8gwDyN9WleNf4BsR
6LuvCkVPq3BEdGImRiIy/YbCkeJ1HSiEdFe9FwweZJNhSX7giIawwN//GVHiKghsl/OllsTug7HB
ZE6378SqDZM1MT3BdZJqASHIHl/REqN9scCS/4TKyG0HRzYig4mQhMQE1EYr9vP0Fq+OWCz+P0cz
jAh1XIcKXjxekbiAc1uYeZKupoMJHIHDcJK+3V7+jhBR5Z7dwhrzW2SIOEeQzn0oU/LFFmD7u+x8
WeDVpypONzReQ6w/6D+v18+FZvCr3M/h5XNeK+ICByo71m3U+njNKP4p7bJaUfc6BxWDBP9t7qtl
ZuYBPlbMYPa29ZwKvBepntL2FBymdhfPSJyytCrrYFsEPHbI3wtzbOaU9Wrm2xV7vY9W9Fi+HETb
1lG68pvi03sDqQSoiS7vBwZ/9iwtOBmnyH4VO6g/WupSj33kulELW9LL3eMQq5DYOqImdhiun2Fm
IGjJrS9gd1evwYfuGHTZkPT5RES3jp3oBhyOP5mVp9ge1wPWEOxXFTZoRXiW3zBs32UBYTWIxNx6
hYhI1SsIBM9n7tQXzJsO+2Y9C8/XVoRPTDNAsi42OIix1MUMKQD3Alivic3m5+hwUpxXtakbJwce
rZubPTrs1q0prLwrweIFwdiM9HauLE4g5ergPfHNJYpj6nwNu1yzh0EZT6t0auXTvYy8P6jkBWnA
NYpsfylH8Eiwkt3TSZ+JbWXMVojJXP0Lyvc/p5WVnzTz/bmaf4jPv73tPxMZwBozdIa1ouTEPROE
eBtS8pdAe1Upwo0r6JGjpaCZXB1JXcpLU2lRJyQOFRFCO2QqvoE9fRO/lGt7Qaq8Ly+pByTNZd4E
yY0Z4ZqUL13p1Y66chwMzuQgY6tMLsEBQGSzzFwfGCGecPWkm5iJ2T8jOmdAscdUICuBkTFqtGtX
bqemhzYgdTKDbz8yt9ZKQ89sr2/F91H95wjZiFgT9/GsXDMJNDw95OgRdFkxURIUZiccTWhN57/y
cqNnHVHJTiFw6InjbdW//9V7fc9Xo4M+bqXUwZoSLcVNWLTCSjZg/6fDt7z4rJlbCdIVcF0owQDi
rBFX/e8x08yUNt5w9W/C/rMIh7u5haHec+aN67BzmgMMRa0HwDhKwROUm1WXgpgvJZL2ph0H2EQ+
YVLSosai9H2d4SuZ4ilpRrOoUzUWsrlR7zOvflhP12MFzC+RnrR9xDx/ViiTEZxQu2673idoYN7E
+4WizJJhWMfbzCJwuMtY8JS4yJN7bo1P6XbdQYoxMNttaORCLsmB3smdOMv+4ZmqfSnC/dHXjhSm
abVIzsnbRaeFXe5uNTBr4LpZlA4uu4qCQHa3b1Gq5aLMKFzzSlIZA+TMioF4y5qptA/i4mMssEoF
FFpT27BUkwujB3yJKQNoVszJXxs2ypY1Tvki1x2BgdWm4bU65q7yQES2Cl5+PrbxdJAVT3uF9kPI
LyNTZjTNkPOy1HQxH8EztFMzQFViw94iigdWlBpAntb+OtfjGInlBHiPN7zXHRHwjrkzZyQ3SfuR
6OIQH7ErHAiMmFBQKTgg0VjGE0tWoM5Tjb8cvTqydi7DWZj6sNmIq+Z1DnNDoNFMbb0suF5Nw5vd
VHkHiby95/mVGNDectTHNIKlDLh8AV7TDvURxqKevyjISNDr1d3ccaISCPUtFZA0jYzv41G+sys3
feTV9LWtUV2E+X2mdf6SBo3ZMgdQr1qj81+4hmaPeLqT/HxYebvqGvo3IdLbgrD22ToYmpM9FT/M
WSCiLOi7JGCT47cDLZMWd5Le6qcKm/GKLvvzE5CDzc/rJ2hj+6dJFs2DagRoIRAt7LO6nFLTR/6P
XGO2Q6/s1zQiVFBFxfBv7wrx7pQAUiH/OJEBC2IW4+ciWRfjWf3jCywxEW1SUbNfUmEw4DSIqhRn
+AKTFFQjSAoFE4KG4LbdUm3Nunnh6ACiqrusSDjDBws0fZqDbuoAOxZgxjq2IzL9mgWe5Z1PKm7X
eVTurjNGK8cJRP42iEhDGzK/0ccxKAS+dagQuDNv5NNiES7sv8CS1bZZ8HysY/61XNIS/dgnx0uK
OFIscCi7G6N9kkxAS0rMDI3GHc98Seyw4FeWMGQIY4Bd9MxxZaLrbLcsshY9NGvN5HCCehoxARZj
GKq4BYVU3tdpnPDi+WcXJqCcQa7PNFPM/GH6gU1r/3JwmU6o9RZf2pBxc6dzz763Djp+HrhuqC16
Ysolrx2CSpc0+XZaaBBhOrBPNOSpXkTGTrv/KupQOZYbTeeNDt7f06HKOMKjNFf6LdRSVc5tKrX1
B2WxjBb9FZOfvL1BDOK4PVSjb7Qr+k824R0pCu3Luu7LHzjKoiXedHHUE4YIdMvHsFjAKhb/AUKu
MwqdAxXdfAbOvtFHlly0Pwd4/rYM/BeZNnbUeKpLJ/55PnPr6d471xWdfEzhvUWG1CHMFqw9BGUh
aSvnjHjmmWk7RgjcRbgKhnFd5x+enjriPSw9Z2yB7WFvAqgdK0wEylOaqlmBDRwcB5LH88P4CLfP
x2VrvqORhKoO92OqoiOXfEzbhFdCcRkP73VyuLf2k1iM8fHdLv9XnnSoHLgtcFtH4xoOcI5g2HMv
s9Gh3HxX0N6eaCZxK3kI419WJ0w4D84p1dDZHadYamfQZf9VeZYHQA0ZMwMObUWGTdXA4H5SU4Nx
19OlnFZ5CJTYD4eR5OzQyzclUqUddj3EbPmD8Uq/LO2u5Nt0hMOWR3LfGypaJPMvgRdtotjpWbsG
fyM6Wptrpl3eUTByvdqwtjyfAu7Ygi1LdTO1ichrVgcCTbA8/Ql2CxKdTCh3SBp/x6dxmTbqrBDa
xjP1xp8VagfZ/PjxXT1Q5B1L/QSbptUZJgo8z2BzQlBJDqs6EpJPdITL/vzxdfwVGx8/ZcccgiCo
OHvC/BPkcP0SHzKyX97nrsDE7iM+vagBwCA3QSaSzlYY7IamnhGXlIUmGQjX5ujt+f0zqkU0J7It
bA9EIO9zFpTmx22WtU79WIqI8kz1+MMwHAUFKBtwvXpc54BXdcweCHBBm8K6xw+UZWAhlttzBWHm
E1LPuHs7rxNnL1sshEoFumm5nI7s/lK0TeCK2bbEACG91y7TJne2L3c8v4CDlPP9bHv3YumHQiuU
t2wTGmjLiwR1O/evyB0iKPj19zI0YA4/QqwijutZBQo3zEARlFy+6HzPR0eqO3VQrx96i0nXdRjz
eI0ZGG8Vxwz54njY074OA0I2ZK7n6C8uh6cf9eNw/uSVBLOLET52IN5CuK5H3ufb1sU8m9ha4qou
QaNtV16AaprXHkBUQ3A0VQtyD8dJ2QYfy4XE1ICjkjPAvHdyEi++HhCKGQB/LZE0ZYRa6Aat0ndk
YwjlzUJpGiwUAqzYHlxf5aPhRKicUQq389AlSzzDum+gFqzapyeckcozdtO0gLy1KoxLuln2pZuc
X89znxAs66QvxcgXw7050mal1Fk6iCTrwy61O3ltz866MLempII1XarT6BsJOLiBDKgnGSs+f1up
Y49pa6X8v4bbKTix/1GilpNYzV7D+sfkbQ5LTpMj56k7JL7ZC4Lfdhsr88ebxn2J3fLIXU1nqTrq
e0SQkJmcYvIAoxNGWAnPF3TROdgMRfDnLMXZgXmebccu+V1gGLb2C3bGIrI3vvjDH8u+0d/7CdSM
GyP6qgPZnVkzl097nEey6wtU6b61rj0OX1ph+OgFeH0GM4Mqi5YOhwIjfeH9UDsgiOt38Sxu8kSA
CpJ52b4iP7uDsxX8el9l2gKHMlthQsJWPnBYDTPqiPIrpTpJNNR4HwlgUSPAcuZD5CmyFKMjZg+/
qnKdbQzbvAFld9ZNc2rmnVpLZ2jn94csDSiJHcSASkH5PcBKb2oug1PGHROiFGeorI0W42niqErz
pwA5PJ+K9ZrjkE3zpZzC0jp12VKcJ7zqfsyd8Xy4Bsirvus/QhySzi5NNefFzGL98DWaH89lw9Qz
72oMKr/ihPe5oioSOg+cCrGxr18ya4OIlRg9xjPg0u40kTd/I7Qy5iw12yhxSafXcxB09ZJZ8lnV
icwparWJeAM6IKBE8HsAl7Ffq+/T6X88N5JHM86qvxHv83P8E54NLex6zs9fpNOnDRtNjKDBtCdo
wsLmNaMBTdhqGm60WVVDHCNe07qk8bpCnAeVkXJSSIqO35M2jfYddUHZ3rcqx6s/XQMkz7tFWwJv
UXTLHi4IS9LWRmkK3fPlOyB1nd7PeVfxOyR9kaaCYh5mAYMLkW1KVZLte2hTCWzzfVPriaLLeoww
qb8aIE9w4ch0B7ETjxjn5ewQhwEMtuCh9/hYhiKoeCnolJvONNIi1cwDklcx/txbvoW3ugwJRWu3
4WIelNdSFnp/8CCp8hCiadzh0Gfb3acCSnCt3T0750rF1AoxXswPu6idNF/IgZYgvRqdAltOIomi
1shtcbaRegvcGqu4BniT+rl6bAhjiV/aiyg9rnj81CD5XgL09foELd3KxW1nIe5ZPoq4BG7tM7yw
go4TPXp8Sw5Z8sknmMQLbrItVrvGChNRb14Ty4QNdfcL84G1vsSaSJPZoT0teFEiK6rYYayuwJ8b
Vsi/BQutaAyQA/unhMMxmZl5TKedU8FZVTyjC0yib/RSFzwUI1NZ64IC5t33MqmGMxLML4kZYQky
4AovpIZpu+NCnBcrjoHE+MaW0HUh4Ng8P17Mo8pFCmzftu0XaiGWP5TptDhDSLLOAbt/9Ld16q84
89U8CuQv0ITYKlOYW1pf44MxCAMlO8vMDU0lHLEe+Oyk+iHePQkYKye8gbP3/O3YRRt5cyBUDjNU
c+s7HoOddG6O6w9lc3COeDO0NljhJQk1ouIn7VE0XLcgiTROGUM1tDtn7kKXQcMW+lUAaMQCxDSO
AdX2EKYbq5hUFbzPY2goHkPP8Sdqer6+Alsw25+gFbQ2ntIC7JZxNo4wYch1LEGtZZxR5VhONt4P
N6rVR4TrRQE2u9oSVHcXxjoqdjFuL/phX3+6fIyNWzgUqT1GJa2FlL76GEEyIfNXt1e5seUDnC9+
c9ikT7I9XQ0hbl13nUyHbbolTAxiKdVI6+HyoWX/flECh249P9MLuYWTveV9eMcwEPelPr26G+k2
C4du+rRJzS5lJC7HwVokNGQbxCo7otDtNc7hgKrbrjzEZ56eGKr7ThonrytK1kmu4ucGgkUd5mdB
6ieZMnGoO5eVx1J+77uT+r66KRTmfn9HiGS2M+3RFY6Y1ZiIfAQHr5dHn7EY8wFHj8KOn8R6vpYS
hui9DUI/9nUjTH88RuHl9Ahc/jpeU0N6pu+9V5el+bJrGQLG7IvhgQTeBVDpSLQs8YU0Wb/i3VAP
mkTz5U+mvyHYwRhdQHKU1YFh9IdZ66+kCR9aaj8dX9dk+7BLJgptzURdlvZqu67qvBTm3T+EK7Zs
o0EvTCLFMfXDg8v1QpeejmgRsjgyzCM0wHxUm2WK2lLOfcQ38noGG3hHTSAGWcm/AMk41wrzksJy
+mi6zJMYBlPzZlEKSd3gzliV820W5Wh+dY5B/qjwyglkREjmv3rfOrZZNNVK4E0p/EYfO47A0SZy
O275W+DJSMpjm6jvqkusaxQ30SuKFmw/UC5HnED7TWSvDCc3dwuw8dnoRGsN2WmgCpZ6yka/nn6I
Kbgl8qWUnqa57jLOdaROMft5sQfAxAprxF5naEwVLAxv+2AbHgOA3ApA3IyAlOsGNhpa9TwU1RFy
bDDab7KqspZkhXt2sTBIyhmHC6srwnCV2UcBR2IfIxQ4lRDu10VUZjbulIzdFMu8Akj4whXbjoUz
e5EIo47okxlKSD7VA+zwdfhlwkQYlwcuvKXSRxAW6x4aqkH2tJOwVGfMzRT00yg6z41e92Tj+NWC
/8k0GB/PTN6PevMO3r2yUy4xrXvENJA2prI3j2y/cjFxBb33if9JvMkp7l4orVLbu/b4XxFcN5Wz
4gr9kn4ynMqMPY5dfeK/3O7oUZGbbBqx6V/ZiNSAF64qJpd5wte1s7zbRWC/CgkWZ5uEdsfnd+Mq
SciT247QOh6MhTmknVXnzagU+HS5aIQzrPlFtvy+SNiZg3iXltFrXiLv1ZeksYrTbSazBqScUhJm
EbRXpd4kOnVL/ZagoMOHntCiucnqQ6pKNvmja9k9RINwnHKvbfrLF5KSOVAzn5ZYNCHZV2NQa1I2
Tp8Lzu4BNmainpj59i9cW6UafmIlekW8QnY/Hpje93tiFDt/zj1BipU1nA19gWNHJ+AC0U+hnwSo
1F3FOPnBzvC/dsIKifkvo+vx1l/n7lpInCuBhwxNnvgImbnzYrvHWHLbP1WUPJmzKyGEYMJRrOug
7JOXlGYpOSfvrwOdynQhM/fRceoZdUPf3vPXD4rDGR+zxmpay0e8ZERrDGXYA/5mD7qy3SDqJXse
3v40GxkJ8auEcQoZxca8XOLgZ76seOrjqqC0iDjyFssi4JPaM4whOjhotw12FEFVzSFaO1Sih7j5
X4lt0wR0K3dVObja6w++AU3iDRpabzOshHHdYfPp2XMikKO2hmR5j7m9X+V2pIGwGA3hZUtXFCp+
wtSweG1QoQkb4P0BVo9dYE6bS7aQ29KTvuBQaGGcJgYlLur3VA7SX7afPSKn1DcvGJrfq9fwPdfA
+z3/AW9CNRaRCQ/9LeZ6AIBSreCq42w8Jq+z63pOTqkLwKmqQ/4cKtCBkg0vyvikWDUCTlMwL3LX
00os0bzs3o+N4GxU/A5yG2IvuFodTtytcdbDd6vmVwTuOtSMuWa0155LwM8Mvt4bFJge9oQzmHVC
Bendtna/VSNavybEjUSxbhNDIzamkopULDm+eRntggYH9JJ4PtfSrktQKyeGH1tnzE+hnlg7XBxM
QXuUhoHQBSKh/yvRVN8DBuXMpOse9OAG2odkFYMvVKRQ1nzNcLX/C/Qclh1ApSdlYVqCbg+tZgjd
71JbCmsFho8eBcSqONhQiLdFChPmkwnBzLYxqWajPTF6M/6guo1Ha5viwH0z1puBy4KEzl5mpyz9
7hJA9jeZSyI3l57iUvRIKS44Y9LzA/ZyLhPAWZ6S4tnGjtrhye1+mkqjhx4LZ0ZSZe2MavKVSyv1
xmEwICoC+hnr8zOsVqVohad24/C7sfLvyjqcuM5jI/7N+ApuYxYFfkZFGi/S8hJrO+qw7jEEqJMx
iNILqMdiycOCZLY4+1Ou6bTG0JuYnvukKvLT27fnxVD/DKr1/S3UMyBEUAL7/24VhUSK0SvQ3VZM
dSABMFYph22a2fe1jRljzObg9IqPM2rT8LqvVn0h73sdHJWMYlKLT0/iD82QcejqGbyywM5wBbfv
AwpJ2NhxRthLmXZssN56dF3j3DNjCObLnALewDV6T7KBo28lb7k35oPkMjl98Swx/8BqC/CphytU
FwAy1xN5jWPGePHGp/TLEkLGOWZ7tdYy9zVNpFPaCrAzuQN7aUFM1c/nZTTgw/NeAjKGY7MrPFiS
VZbXoZt7p7gtS8ghiYKbFn+7QHGMT9169arUtFuILFuCxzdB21E2ohG02HgRfdoIO1veuV/1Yp6a
sk+A6dWak0yxXma1LwdkOln0qL3ngIJObItA5XcvKAT0gJ4In5fvz8THBBPZTHk2MnCJhFAIjr6q
3ec8rxOPVHS6xtYjvNxqaPmZfVdeuYjBMu1z+moZHfRKExVt+Y0meOTHYOm2ZtJfUOEKVlgYu72V
/kMyYvzDfhUkYgTQ/zCeqAJleHW0KgTNF67RmbWwkAZRD3nD6k032w1//Z7JnlRjkyqrsKpIapLd
BH/qUKkrayfa+T3iGDkBh5Q7NMq6k/+p6lZQDptKv7aXi9/TBge/FBpxYbboMIu+PzLk+GzbNqCk
sXukX3lHh5F7p9rG0O71YSWJBPGOCeGFOR+zdelk4dT375vfHnZfPM4XMzclqjrGsx3ZnewbWN1+
hY1DUmnnSMAS/eZ7PBJy/6sdaI27IKrMlO3gvB86fTnGkXmAxGy3MmSojFFTwDOTIP4TaJ+vcaZW
qSh6ozZHJpV3p5WLmeL2SeSQg6iinFoq9hmxCtNGt70FEX7iciAbC4OC3biHaCwFPbfk6eOfvaGK
FBEA9Nf/h2uSbdLaKzoeHoDFzeS63ToKN4l/dCWrSj72Ag2+YSV24Xxpb/vmN9CzsKiDe+GdKuAy
KK5waKNFIayJVlNQfKOMeZJ853t8MOnCkItgcBpgbTrolEv+jIM4Cq+Is2OD3+91+xC9Xm+jhnVe
chZOKj9sVDQlJHf6QSqefJobZd8F0zMyuw2Tdx3bSoyU2ZeNm+eph2+2fxD/FKyWTEyfmtqc/5dt
z567i+geoMTcDap93WPz4RXaNXn/triB8vehwiXH55wDzW3ZvUAfYPvxY+9iEJwbmacprW3vnYRk
rcJWGCF5DKKIfQvAp0sB6+Pd/vLmFP8bWrjDwVfQu1t09wOqWb1LcuHvyxi3ZdJNerSgFPx23X4p
U4Rh5F1QlHLm/uFhxXrF5Me1IMTJIoMz4jgPV1ZVtpWaitfGyT08Px4asH015RvphiqZnGL52b4y
NPmUoDRbYpSJG4nxfY7Wh7MaJldP4dPJgj1ugaZLJfrXV9zZQsZsVNB+28Xwnm5yeBrtDwG0/VE8
TjBWvDQJkOBvmF+/jt+DnPnwmGmQBcckT3bOcf5LAaW3lGvRSjM8xYEirBGe3rvWstsaNDwOqCiz
FniyIhCHtSslVxOv8SnqpRBDRVuRWSjNsf/eHn+NHc0pHoIDPCqkcGtqPF+v9oJ6iBkCTdSR75ao
goxxbZPjzutQLgJsEROO7FO5wDBVIzT5asrLTnMHF/lqw34jYXyCfswXXAiVSpFC5UB/6Sr7D2Ba
65uN90wOz6ZYoS8cKZ9DMmFMj0S9wlFFeJqTdOOnGGDdESbu8RH3ml15KUTUtUj+Jrg0qOc4d640
x+48IrGVjpqyE1wRCVzwztfA4HJxqHAxxqRdW0NcrfJuGUDD9HGomJek9cWq4rlrVnTIyUcsmTPp
XCvBMxNcp3rhHg/KVHbX4U3IECimuV3FFIXpQZMIDecA9hV83hS4LVRl93uJQwtISgjEp8+5yTNq
O/01MtlS/o6u0FPjqXJj+oxwZAUOQ4xOypfTtrDkrmRn4WSLHB19HDsCAYPPLIkADIpHql+sIfYA
z3Mp9UtssYv3/cst2qbdgdkqU5Q/yDRWdB3gcBmd51k1RL6cfTg3wOT7OLctjx86eYCWoAsBprTg
lZNsI7zlRS5w+YWRZ0XwP4cHRkpnLiFNTc5/+8UZz1O9FhAPUU+JGx4nsuT9yhQHdoMa17/gb3O3
reL86j4i1RyQBpfFCgoJceQCEFPKh3FLeDMN6sADu58LCdzodrYg9dUbo6kinn53cAtsq4QdS+6J
HAhCy/9zxc/RwV3C+HdtfOVQr0npoGpz8fJG9IPTuGhUVVw0OPW60LqGWQ4F29qU34UWrbJdf9up
oNY2b0Foe5YgvKa/YQPdR1jbYKds258dzbvInPhUNYxQpqmJRXS033f/VQQKgkKk6vyfU49KxdXb
znTKt87eREuVbr+6xSJtbouy1nbrJwsLkLnJttObidZDsBkf9GIciFU2kkfC1jgwweR4K+oG0WBv
FUhlFXIx5IKqzzwzoDKuOIM/JemTXx/gzW8TDT+F630WBeP3vNNXlBwAp3rruAY0pEUcgSmJzRVe
VYcJbQ425jmWC1NQK/goMJpslN1N4uLGIfS1GBCUbzOVLYOEykUxgqljdJmCrKLF/uNzX5ZTYPv0
oXTczyBqO8ZECGSEad5qi10QuDireRlEzv+s/YyLiXmVnkY+vuMI3jUk7+v/vI30vTrYogpZ2ws8
p7fMgW7TxeONTo1RBzNc+i50bEd+2uJDaKOiOHQJ0bhoUH4nshidFLHnusSPeM+bD3oams+uhXey
hHFuVMHc3+8Qb+HTVxh+p96rb81lIRUBdnNUpJcDv9XYgN/AEyY2IP/B7rvacSitCD/Aw3y9MWDB
WincCRG/GY09GRziJy5o50i7DczllyZSg1Wi+w6y2f/QwZrveen+nU39gp6raqKLB6qwVHC9LZ1n
sdaFowLZvcwb9IJWuTT9H6+4AV/LmI14vvmf21Y+Cx5VOM6rQ3wlcvycTCGDE+YGGnVMXN+9vFGz
bWfi0/as/rndUhx8siRJQ6VkiuM6sDALg3aUnyDhDPQMPps3IsRGvvwmFCRf7BxU81zbrO9q0kwh
V8HHQi8uvIC7vhbgevzSgjWpWrIy8tVZ9/2fxXvvxe8g7ogZIHdRx+s1Bz5YXT2tD5t42D/uve1I
IyH0Z/siCUtcyZfRETVZFxFZmPAOJy+b1jP25tnXnixfEbgF7q5PGNs6Dt4Y5NW7jHAX+qLz6b99
jilewHO8tVi4U8PcQtW7ivlqoQ3Z0wneCQbH32eEml/hfBmfc6sDjn691n8PQkRWWt5UdR/lhuET
QYTLcDyMWZLUyf7HvfSVudvO+zxGXVhGuG78gxEYbBas4CR7Xj55OPHdw0iHBWPm1qXgof7F848G
ff29ULaLC0fbnMstxnLoUrHSVXJuTn9fzwyp98Gcfa8gKWlJyCKmt5enR+kwTb+UDB3DBvs4bQ3z
BLlsFygULwYHa7oAthp6T62XCMkB4hBQdmLsORz+Ksnyx7bAs5wcLcnc/Ca9sPTAMvw0EWqXM34I
GiS6m2UuueRthw07f9vDCMfGqH0Xhn1+NuReroaLAaen6JLpALEumgE3+nd6LpxGw0Iv+oi9uSTX
EXXalwtqNCAQNMI1j8lydtaHDu/vocXQxq6p5g5NjiHiy6U5zOGoVkF/54yaobmIL9po9Vo10mSu
OcrlqcRVOYEvg/WGocOTrciNWVzopnzK9Ge74yjnenXspUMHHEbWPujLiiCMn3n+PR6hnEvaTnHl
UhShyv1gR4mnasG0nCLcrpHX3OhNkr9STJX+5HrEGy7e18lBINqqMD93RupiBsKAFOZecmYBxYBy
G1K1WGabLtXdrajgGkBnCz9+DHETawLlg3A2JTBi7hmZKv4yrEOuEQ5nLhJZc/IuubWaJ1tntzwj
tKy0AHZWdTjm05D6oGREA4xhs2WhVhxkAqobVz9D56Kt9wibxXAiZH78NXvH8+JFRFuqc4DKZwE5
5tuKwQ2dYW+vbkBlLDF+xJVm7kJSd4tbpZpwefnz9WhSmhRGtVLryhj8moZ26pI5VN3t3c8irZ1w
eUV3VcUoxR8OBS5VjhE5kSLhTY/6pVnq5nchaZ9CoTz+VxirGEQf0B3fVcMoR1g07reKMR6Lpq/C
SzN/O9pFfZcAG9wOHTJmlodDrkySAPvY1GDYYBjwpZMHzMvGl8CtS2IRmTEj6SYe2TfCq0Ahru4S
PPPyZ28bRGNJo58RsyRADDOMFBSwNa3YlsSykKsvJR6kC/SaRsWR0UGZJe0/tnrMIjtuold2dWUO
Q4cKA+cJY1+aTUPjXKIhxIcaEo+eAzW9CG8LLPZpXq7LYzvzr+wOPWGfjxLDx22zbVIYt0meUeit
ixd15gYDyZk4B0iRQnfeCfwv5jkYJpnrjn2Hsrh7TE0F+62bXQeMPVMKFrZslGZD7NjrHp3/kzQe
25MifRtUux+Ht02wC2VSl4Y8OX2B6fBnL6D5gZbvqXwM2ldZnytmX1rCdCuf2Lbd6sH6r+w+/I6e
WWWUEDYkfLlTdEWGqatJkjk3GGAx3TWDRKAXXp4aK8NkwxYcYejew2Or9z3PkCBFVTo5P8x//Boq
zv8Bknwt3CLA0hbpJVhlRLoBNsdP4pe3Fe7QUkWpUQIhUbQi40F5wiAMFqE4iDu9Ml3pnCRLwGyl
xXDcFlzMNIxVxmXcEXG3+4kWFGha/Jdc9fbr/Qj+S6okqVW+GgyMuAyXP2poq6IGtRINN+w/xkBK
xXtW0uEpzEGaRpzi55B7oeQnSBbHMrMhdCltrjfXhFb7G0aGprPd50+Q8U4FVZTvHF1bMWmvAONF
8Piw2wIV2UH3l/OacsKc1SYuWq9CT6tn1bHHMZQsZ2Dc8jsD/S9iN6K3gnPc5tTreidhG4pKqGR2
EaINHz74y4vrH1/y5yeSVZIAJI3855W4ebqJsU6VvRlfNeTGD0/u7CPULingctPJwhA89T82IcWA
wWWsdJ9aKf+5irBvR7RlqGRgK7IZl3+bgs5ZjbNjseyBCxHXuJiSA1gzRXu+bO2z8aI3EgG3G9l6
ulgw30b6SrUOgSXjHLdbtTQeqdUj/DVSoma3EQGnaUVJQtjOS6VUP2p/plUpeazrfgoB2+OnAWHK
esML7XEuubRUNL85alSXHo17HQYKhfnxG0w+eXAxWXyrbxa0PrUAfeqXFgR4vbWCUJkhIn9YlTuX
ZybCA4Uk609XRcj0qG4y5gqcA6xzVU3a2sblg4Zy7NqVA3+xZdpfExN9YgbRtisR2lOSoH914CDG
HwvvihcPG/RRMbZ0/1ZojAVc0+l+QQDmJ+bgl1VkYwAGLcYEgFtIHnLJE2/3ctdaNYbAzvjbmGgc
XjajVw/CJwCH5W0K9x/XCg2Rev/yM3ApWmpamu7nkcT3pzG1P6Z7DFOPJ7vr652nn4D45jT+Cu5y
ZL8PwycEUseWCVlxXXGlQAGeMCRsfqwylrZVnMIeI0Tat7ba6FWfWV5sHHSC6f+7lIKv/tiZp0ve
J3f/S6+0aWHUGAdoYA0CzqeBG01nLV+m3zYXJVgTD3OKYmXw9ilRl8g9npvKC/6FB4dQ3+T+FcN9
YFbpHSq6LdzzwCXyLCEQjCwKoZMcb7uTuwaFziDJPF7C5n6c04pX8QoTsTDr3bvACnr8ctZnuucj
AHKHBSpIYHYq6jK76Yf97at9YzCPyGXTW1LQF19/aIZXyv85CEAvrQqVIA2HRTeGwCfcMnyNb3ku
UBwc3zIQLzkDuaqlcDQlowWfKTenMlK9CbWI8hXBsf3Qb871jTB5SRNwzWIMps9wICHAb6XMBddG
FgBmqn6B56V/evAdr7D+LsdMuwFM8vUzAdW3KhKr2ft5G7AJQL+qwKMM6YmNtEQOpXzqu0U+bRQe
mTCTDb0uyfFqAsBKE1i3jrZLYARuwMU/AOYn5cfcukwXcUiUy5IX711wGTl5Q0GwgpCnTYWaBn/G
cfoBYrpusQbuaUfgbXaBK6cN7ErnrO5jQnpNuigkU9J0sr66FxKYfp2zYcvoV7yhIEcAaLYVFv3T
L3Ypaq/GFtJ2/f3RIL7VFVWMUNSIyGISVyW8VFzwyolHsHnoAkeuzlpRr6BAElbx8JhJQhFaWL2z
NGcvESyOWpmIWL2tBqinVGu6uQuhnc7DxfCWqcXs9gvf3aXCrPZFHpI6Hma/HvUNuZue6iSIwFsl
xUyVfzDg12KAcb+fkiIW0O+MhK/s72o5LDtFRvAF1qgR2xd2//iTA+Bpl56EFOzi3Pa0VHA4Nq2n
Ci7y57DKhRkh9OIHviQJL3W/RPlXK0ljwOWDyUTQ+NZ62R8fihRzYih496JMHMoUDnu8XfQkudEP
Wm5eOap0+oTymSO++a9mZvy2Xi+o9N6xx4dazQjJQ91qYmZ0o5rMGCgkkrPb4DFczb8TZbxKIsiZ
NWLcBImXdu8G8KeW7u4KsMyDZD3pJLVK7XGg9dwqJ7jLTNDFvpJm1xUJI9MF14Xtkb6qE+v6/7/1
Bqj0nJ6eC5jY0wZnqsa5qxNmNNK20JKxn9OysZxd57qnGL7v8q9NkUxnGNOqpHpt+qmzhR44PSs0
jMGGFkAH2ohgj73uadENkXuAOJod/G4CVpJ3bveuDyV/27KFpZmsbB/a0TBLLaqajyX2PrmzFs+z
FoEAOnAdily1q1heKZvdSCpuhHUmpUMbEExtZtujvpKOVm9HbW6/nB9Zg2GWerKGmYUJvamEU4bI
VbonbcRnPYm3QJts7C39XWJvIg4hX2Ft/NjgwjoFpSeCRuhUft8RG15nzm1a9iYk6qhpkQIaneE4
E+A81YlbSlctRtQMbKbPzvh7QeYNyUm1EvWoy1VxuacWkx1cw6sjkNVC1LxghFQGjqb+lbKw0N1N
el2maOiwnK4ZgCWaM94hESdVNJitMrwwtWqKnkHfF9jkNl8OswtNhm+tk4pQYXiH9nnJcYHj5aEw
xund8GE3AuTk4WQ/tQQQ/IcBtl7GhXuDw7q10bN7/c1DXksHhh1aU/pK0llxo0bLuyY0O85/w3jX
04/GGunDimvpSwx/tJqJ0YJ3JErJwXIjpCCls+P2htSL2xy64l6qIJaK5jvzbHsFhKrlpgStYhDj
YnYLtc5cZxM1zWZaURO01X1jo8MsRNnAROxl1gAxmQ8r3X7VgoflB8BTD7PUcv+XASIeuJKfa6EA
l8yHaoFRbpGcVqG1l5AzoofqKMV2g43Ejmo4C09G9G2GBxq+4IN9JfVYZaFb8iUidwaDJ+HhhuHb
+hrJE2gTEBWTEU1/OTiZufwZwxjG81rVaF6BUT4t6Ye7eFLadRv8WQJ5wRZ2dbPhhMpL3th0LIC5
hkWU1WNjOa7O3H5EjUwAgpfzaNr6LmfdF5uoOt7oj6I2h4CGAkKftia9i6GiVSLnYhMlznc1pCVa
e2gF+ZEPshh18duA74oHxZly5ygt0XiAmWdP9wEAiaHkxUPgJzNkDpjFOYA3ld8hfJ8+Sb3tzN46
vKf/Lp0QWKd9FO01q0kUnraM/iAq1P6jVKIURSSzQZeQYmFkAa7GLdtgKXwf2tm0+QXsRH2yzmpf
CZnCDT77srEGuLlnpR/hr6kfp0/5XJl813VZwa0MHbrUarfMaeRSpoaWTwcqRFqe152rVHJ/VkCP
g3G7CHU19K8z/acz3DfytMIFaY1pOqOSOF8dnv67IDq6dkWF1nHe8scdUW5lhOpmfW4kBoy8Lvyr
np/acyMeEhi5O65PDFyYyTgJUhYfoAn0Ht4kJhKL8YgaZmBsFrbCJE1ji+EqwbuGmSFG4RHl9rFL
RVZJU7siPRVff/ZJUnpGIYvCNcyWkGxDKxlyChWPjYpRON1LKq1AKPF6AXxEqpViIVDil5wiiAmJ
v+zoOXJ/cDfzlslc1yWBpuXc09p6W8jQDy7UAIT2fSzXKlkunpvxLpPltCWjfBVADQoxLb8CJPij
2HT0eG0D5Am3/JP+VXdWNvpfPw7bCOUBOz8Ynff2FF/Usi/E5EWBdvezhfGqo0ydvBvEN/S32fav
lCApnHxQk4clHzngzY7BlDJTlWm4hdwqfarOH1VhjzxiGZRzHmM/RxdevzOKSAvs71LGvLYFYYfs
9menHIS/RIra5r6ZdVnCdMNOEqx8ObFfKE9Ww793XvQJJeSwUDndWXCgWwxYBrKJ0q4oyiqtpv8q
7dC4mPvT8xALFOIw1WX60bAG4kRbKJHmmL52dNSyzw3pQ9sscODPNFv3QrbLPu7/VM7qgB/TMhe1
lRoY2cSj9QmSjSVDhWhlRXLpKD009rzM8Cxhz1MgQihRDKs0RaDIQMQg2qBSsEjluSLI/FwKP9s4
uOeU0dwSvTValsFtoutalT9puwb+5JI3HbD+wij4Omv2CvJhslAt91E4/CNbZN57mZoEws310tJj
tvxbJiEwmqgQreD8CBPbJ1Vaom9hs67qmUv0s/o+mMDRkDfmbJyHJVBYVO7jQZzrmhMXGcLw6nud
FbGxGsICMYoGyE64uq7ePhnJ/i/jjNB0GHhsL+2WFvWjWBeYm89PoXfehZMyd6dvQ1ZOMhftcnP8
GFGDg8qyc9GzH7GuDiW46+B9AOZ3Gn1XKNzlELwjiP4feOr1zkIUzYlkJ5JHDImr2DLzIpGcBQrC
0P/+vTS89FypCNLsCYy5nZYOQeMSlBi/Oo5+4HOGzexQMeRADiCMmPyBnuKHnCDL+1oxpj6JVh5O
1yfenxCerMtZ1ImGIq5RGpSMz8Bco3tGvlitmWbLN+6nQGBAeptrtWGUpDZNS69PftRR1mKvP3lc
f6Bapu01VsDmHwXfDBr6O43O+qHELO0e2SJdUrs2tf03fnDV5JAajy5Rjk/GnMSvb5LqKXF5jnN1
1nqyX0Pd2G4KBOKJ7N7DzhaKVajOZh2xxlvmmAjP5kMFGMnHBAIubE7yBmbkU2ASOgOR8kGTCzC5
88H/+67QdKFZxHqYeathVHSp+M6crJYeQfkgF5XjJV9+bUPt9TY+D8WOPWVvW7e3XOXGNQMGk2zT
attqtd/aBRfWWMwzLTtMsIyT4fICuYadCx6l4Vzo/t5Kmr79DTqZr+RTMP8HHlyMbn8AKMhCxk+C
JweY9XJylnQglFK1dRoPwQQHSuJmtnOt7LmirUWmHxEKSeW52M4pN1may4cJJzTA8zqfkJF3VyNx
/qIweskI5H2htVuyTXYvkJGYw7EruszNBmzWkSnTwXPc4SDqyDGgcTjf5OrV751FoupwvnsPzBHk
RU84z0bOlpS4L8kVOBD+CxDkxX+qBke7E9JMsVK1WOriS+ENvZW8eTAZiEx1RKemWnblXjqWyfUP
hAOrjXvxFuSnqaEF5Sja3kmUhG4F0G9ZL7wAJWe9kdcuqF3e7SbybxlOtHuQPFcvpSSBV0vqv29a
nHcxAfnoZfaAIxy0mGDmk9xeYig4tOD3RaCkN1TYSfnCF7yQsm9BSjo99FgeHGiiUdDzwyZd9mQP
FMSjfB6KLKVKhfVDlzs5PYnXIiO8HDu67pWOjp4GFWQNRY63+p/jOFpNgFurlDZQ5hXjPx4Er1B1
B/gxfc5jhrsSMbGkUcalhbaL/Ij5BwHKdwh+dEkIBLzKcOsUXkPz+FOgV6Nk4tvqtNDtZ4t1BX3Y
1AAb6sDJcWZOAWfLycVsO1tO5ntnTqNfs9JH3a/CG2uyyF1G1pk5oGrenXop1hmVy085Q4bXnUml
XCvjsU4vNyyEV7JcVOGPXkl0BF/H+0iBDbyNO6jVf65ITt0eBKKCcO5+84DYJVUVzWvy2OwuwiqU
F1YHCulib7mIl854bpFyjSE94DEEZfbWS9R7XdAbdYFIrJtctGx1TGCrG4b3pPx/gvPMRV3mKbDf
n5eQFX5vcnjwGwncNreImwDi2vs3qXG7Suw/4kbj+U8TQVKAZoseTwXD4yjwFeWfjxPSrLVtHHnJ
Nwu5JETKDC0bhUfBGVaTDBHl0qs/T/OXw5vToDBgPq/O82hYfpfTHIcwu9HhU3YmgEibXpon85qK
D3lFXR3YXwlFmwbruMqIeQGqas8TVuygviCxbDaxIi7MkcauQIIt4ICCp44ou33ByQ1yUfIcHgeY
PB8KWYaDz9iFAyUsa0/FQRegwjPxhoh9Qn4mEnmSYdQK8s2VsM1RCXE7is0fAkWlPPovnUTP2/UH
/YIugUwBl3ha5IjWr6lMVkauAd2z7GZPrOvGaGofbOQvW+Cqe5SVmrVeJNjm1oLpxR2gkXaR+UQg
BwiCm0g7cgiZL5+6k8LE5fgC4VnlI7+OOAScNNCc3FBJwR6b18ApNFQbR4GvAeu/bzXUz1LKnxh8
nGGb+i1NTzhVLXAjevtGM42uY9hKG+c+IAuXCtCY5+tgo2jTTYzlcN7e2Lc4AEi+Zo+hioGxoNtC
h+fVw7q1JCqfXNxq4sjqe8tAhUWUE1S70n3PTQelx5qgJ2eQjOBiHbg/2Y4wg86y7CJbzDtvmmXU
qCy+SIUGFT2Px/2zjnmLX4vbMFkhC2wMV0auaWtiZS+kNfS7PTY+ZdiwuiqupprDZ2M3oOryCR7z
TRA5e9uGIGn89B2X6Vsg9OFhM2pdnum4oJB96ITLvPOaeXIuiEWOOMmuPaFZrPAfIgy3WaBf6YmY
s15DDrElHE3d88ZjLNUzAosXl9PxVaKTYn+tE8MfM9kJU2aqBCmMIQDP0gSb+AFHOT6zluquk8gj
NdqISVIGjcR3kDcQJn8cR0GyxdRI/MGkk5p2qH7l0sPGKGQsjm0TDO8sK5upU8wv4nSn8GaGFDA0
6y6xS1iTbnZG6ds7Qocqfol+WvZwDthgueC1+7I3FmsDUl8kyimiygLNUkR9Mky0d9dvGJc0EZMP
eOxuAtd8PK0+xPE5LPdQLpM929snYE7kNbridyWZ7irjgCCkN3/RhRfSDXLTmhfyEf8fpsj4YQh+
uTW4XcxsQvL66lbOVrT7JutLRrXBeIca6gAJcPccO8Q6mkgX3Kswp+sg3rO0QtSpMERsRPhKkXAp
n3iABrwp0l00n7IWLMj0rfEZX/Cr3oJIcmIMhzNQsOQpOOfllxqeOAfxsIlSLrbxt8oU1KNtmvNz
YDML0mFYKvblJQYTSs+9TvMJapIZAmKB3jN60mUCPVm3EytrBWoJ6NQ8THXk9FaDqQTKbUCpJNl8
0oHB4erNYXoq1fiaD5BHx1BbeQYT9JbqolXO0O6cJ0ys7ItqhZVWFVIoXBANATHxKRQWH1QPqIpb
vgvzy4uJY/ELOmLQazX1u3ZpEcCF7RxyAmUfl0qcWVfF/pWqgtBXd69lcBWJyNlDncb7U8++lj7D
kfYf+x8YfkcPyANhv6uuKTxVqVuKaVixL/UTExWAvfGdKZfSjFjM7gvAjNGt4j/fSm2wtJJMvxbT
zgKpdeSDC4BrMDi5XDpgPBbUtpaFaR33rloP4TfrR0KZEOQJSHpsVsKLaMdFD4zOVBdt0ZvfbX5v
zFj+E2l+3FtLCibUugKMbH+56GVX4VisrpTyz6XcyUftspDk0bku/E3uDvpnJ3qtsA1Ho/t4Zej8
GJGpGCeuEXRn4L7iCmxl/HK1JBVYDwrKg6E23i2dp0ZI6zQUP3ckp31X0bNbYkySYt+o88itfXqB
JI/VE0HvOTTOoeRbubgr8sqe3QM+X+GDfeDVz3QtsKu0+Jk9uvs+R/ki6RYOWfarXdQrC4y5J9x6
hD0RP+4yGT8DTKNgGJXZzpKZZi2Z1HGuYon6aRUBGDSoWvyYM2AVTER9nolntE5K/ZltlhotF5/8
bjjir8gtByMnLwdF4sIzfpqeiZBTlT4T2/zbGDpnn/tyJ9XGYRCyZsMbxMi/5uyMgO/sGpcHbXI1
lbYXLE66zLB3pfGZ37kRZvq/RQiSMEWzUAeaif08iG+2ktFY+meke0EUyg7LxEeQ4Ew90Tq7lk2G
hfLh6X32iupgPUARKqYNg3o5u9lKueb0LYGXpAaXLVuX7xVwGmKRZc422FYsrhqqKf3ckSKTVSkJ
Ry4G5ipIT7Wyv5xyrVeDa8frZZQ6Dlom7HrdzY+TBdsP3Fxdr+tNeNonQed/z7qN9ulx52Ujd5AZ
jJcLYMumuxYghoaMvygCHg4BV1fiYkLU7h80c0pRIhiw92xJf9+z0WEGJeTkalfcryWmmblMm5VX
234YVbv0RXGkSMcfJcXD4khwIMwRVf0omIA33sqXkiUFtI3/FLSWsy20HKQGNQl2DDQLabfuXhaf
kNLLcTmD4yN8y0daXwV94YYZ3BAfsL1Fm9sGOWMGvK5O9Pu6S+hTZzNZtDTje9tmZrxp76jcaV8T
DAL16oOUgImQo6WAPTDRI+Q9yACRnBKMy+IIgXnWQmhXL1qXWKHQC9mWbbcsLhJvH08K58xjkkJ9
dNVSFc2kzrvnuzFhVJ5VNNDAyCM9t/QV3n9+O6ai8GBbYvfvLgAhRubDpOciCX3Ew3gFK7ts7+gk
wcrjhBSgmkjtAGuZ07VgYaEcnr3a0kGGEVMvtUcTVHQMHbFikZZPEKz7Whcp8Gqdo5r7/inct6ad
P5nI/CtGb8M3u80sCiNViT0lJOT//E7MV4ISk1eLc2MCW30BKNrLsHJov7g7dbc9rvd6mzXcHYdE
kMkMEKGJYHCXRZPJB2hdZBu+gjuZ8VmVHzrLMY1rJKoLTU7+uWTyaCyifpGp3DKsnj2MH98t1PeG
xqXCJhwtpmRIl2I+zphnWE97W+YFiQVZHuL3BV2Gfos7MlZ4NTnuFWCNkA2tLp1BsnpfmlwAW780
niR7VGfWGJO+UC8NbUITQMCImWWZUDdqepoa1hdI1sQsuC9ClZqdgykywoCg6XJhc+hwmhMoWKlB
KTLwaYww3uISFpphEXq0GyboS+w2hOgxi3Kovo2v8ZGV74zt8Za8G3Z4zk6wx7dVrjebN2KqHXIV
SdhN3hv/kAYKqh0nZoNdQxPFxQsj9VXSI87jJlTKFHYXxUQEJWOeSaUzUw4fqIQpJU4GprILEZ52
JjDqnsWz11JiPTZo2OKOvre3WufpeF/OusbsA6s+aENTEmd2Df5agWrucR7cnccnMlsHapVFMckb
MrSWLlME+hD1qw6CBHPxLxffTlzNjHmUPEaFdUQIyBS6eQmVX8cW+KbxHJmyJ/eXEo6yGaToWQDa
WS7Duff2RwSifhKMFIYVfndt4KcBpGYk0pYAAW98yVv2ZvOQqTF0WLRZMM0cJE3e46Q5rlmr4fNO
ZF2jNtgYkq3+p3r98t1ga140Or6qqJRW05rScPhumyBJONBkDmJsgGNA5qHiAkokY5frQwrVpois
pr9Kza3auSHdQ54Y1XWZT7acKZKS7xpmQY5yNIa7RnQHjvhtQefY/bWo3u5ALXkatlh0qQ5MzXuo
7kn42XQ1SAvhk1dYosKV49MRa7nC1iRL4a56U8QBpYgzcm+3qrMlJ1+yd/RRqbklhaKTQ24hLIYh
jiaxsHWQAfHXRx07YPhec2ESlFs5H7oDkVi5RTfInQn7dHvarZxlbpBO24LF14+F7Ou1KYDN5TeF
szZtHFU+O4fREEJYofY9ARrxBkIRgxhXHhGov9Z9QGGAGb4aYxqYDnvwAQ0cQbSMsoGDNp/wScT1
VN1znDmxJxkECIVHg0ZJJTR8fwX8UuMQRxvPoupZ9ZvNZ9V2lHildRvaqOpPUJqVCMQwLONu0WVd
4DBklTJ+6zuRa/fEmJJDb9+r49VmXWpSxsP6o2JmvJvs1ufDe2tqYI8us1ZKawnN+/s9xmMSsjsr
dItHFV4DwN5QEHEJS6f5Y8j3ZglD2wHnSJkBKi2omFt/77gnYgsWaqNI2aVR8qpvIAb/EGTTEsbp
eTfrZCdlv4FsDIIy+uFQsGQYGoEyceayZyOhhBbSwYrhHUqwRsEC3aPLrC5MRJrtHKQKfsNwGM/S
wsbImV7diDfyAXO4BylR1QHTBCNJnvmCv9f2GmS1yxFZc9oth1c+2Gjmoxt8HHKMqGQ/P7hP/kxM
J6EApMPkdfAkdmqg4L5hD80iLHZy4im4dsFeNFglNwqFPX71fh6KNOSKjP2RI3AnFbLrmcQ/25+w
cRFmgHevVS7sM562y2/qWh7EVgJZo2znSomBi2S0AOjyDPRzWK5HhrsSDOO1hPtBUiWdSyhJ/4xr
d45+dOOmpjWK4XXuwvAs9xJWpmMb1Ma2plKrbJGiMY9WxYKON0FAnV5vJIVwNJgQpdEA+eSeD1VE
GVh75ZNe29g4fTM5HclyxqyLsw9z43KYRh1jbNQgLszNzfgdn9rR6T5JSjyRMbwIwyFDau/HUk9v
BVE9Wb1NrByHVVCs1E02rdZV8mmBrM0mER1y77sejjWwElfbXReDh2xTxXLDTZc5azvbOnuCnKNJ
RZmOmKYefJztl/ynu0buSw0Jvv3yH4rHoGtu3sEI7U8XcV7OY9LsaJLBn4aZsCG/0WNDq3kkVIxd
BqF27e+/QVmGBXZ9XnbCgOiqJ3WY+layqp/b2OC4x+/otBOYapq4aQ73Y2wCjUDtV3DaER+hws4R
oH3B/zRitDK3Oos0gduyzXaQ+WyXxqHEkhGSMztO8i9sADJybJwO3qBVUlHW6XvQcZahlvLRd11z
OX9W6XzJcAHWEEPbGmnw7GNjtR8loQpejn9gvizp7P+RfKDSQSrlxhw96iEXQiSMgMo5Xn9ltbyQ
CMyUleHS0z3XaezVcIu6J570hUkFIW5AgqyetNzY9ZqkLr7CVKFlgAkYD6OM1G2Uk/gyPPO/Nsv3
r3IfwRD6zzqxsZJc6Enhq1FpNRM8/4HrHT2Uqs0LgM5RNIakKbFZ+RZxo8RgmOhRUQ7mGDNjhr35
XXmshHStzDrLjy4TFa7XS+mAFCkhWjHU71lu08lTwke47REgdswic2xuW4b/CT6W99RjqZrqsUbI
eEc0BtKwBVUgyBHu7h/cVjr8shX17tBnkIVVPnPyJPzib607BLgasNjB9zfNPxczIxpgeb4KBAh9
P+NOzvjQm79JpKNuIkcguGbdljkwUMsVGX3wxtQYpUG4gGBg+zY5RXa9c/CiBhDMsSJapsCWcLQG
Xln3tlxR7agYz2GsFru4DmS8f7p0LfFUugdHyl5KI4AjKHUGH6H0AG8jZJd8Pzj2iLYIl1jnpCnE
oENCVpdIOQisNxEzIuAmIAnpd01f/LQxZy2WA/S1eL/z/VaiXwtZX6aKAmtljqh9dnuXy5LIKpKJ
Q4GkyFNMi4XWVoRu1Dht3Qy5IhQ93AMGLBhgt+rlKBerNmBCj1a30ElVS7TMC6aJWLG1JHgq6lHe
zsbcRiSp7RJQIGsIG3ue3jgYkqWHiXpX9SPCXxim3Leo3RkAe8GZXcabE7neRsjbrn7tGtQ3A9aF
99rT8iYy/MrPtj2ERyYaPKKKrwq5WALbp9WVB6TdiEKhud99T90HwbPg5MWSHuukwxImbXQhV7do
fVk2YcIL0GpqWFySBe42CxWodhGi/tlFoaSBey5z2Ty2Idf5RQb7nAlJW48QicQJGR5ACamNPOAw
77hsrupXJLFgPJbsLFsG6SpImucInntk9F/qM5x6BE7jPJ1DSZVLO3mdFcshHFjCMeEShXq0OAYK
Fd8FnUq7UknPF5a84HE8fFMI+TjEAf0gcA1/LjJ9XwuR4d7BjK1ZsAUSmBAe8UytuvuJepZWizX0
g7AD/JaHHSSBEbH3Jk6LtzltKzu+0TbSPPiiGva+rs/IXG2EUTjt410pp7WAcZTZI6GcFBpjAYpP
tjAKFXOzeV35h1U5Tmkp6pAA3paGk+VisEZS0MukkpW8xol/LfUu0eR1hPgYb8nH7+uhBZYvUPS+
aQJot0OBGQ3ZeI62k9eJYC4qnLgHkzcO2A594jCJOT7qwIsDUrFCzssMTVCL40c5XIL8lqoTHrbk
kM5mMNpaX52YzsHGlqKu5PyG5oprRUpe7FvgudCxkQYGLvfnrjtbxCaH6L/kCKV4zUA89k8ud4aA
0+n2ya7w/5fdl7olmNk770kTgDvDxFhTRRKxFUgOE5h5LUxcblRndu40nGTf4tfSkD+iNNdoEIw7
i5BgUBueimspHpLAE5TWGi6dPuQqo8Wd9KftEPTR2NTEFRl62ESrU60KxZphCbYjyMMm3ON5QWs/
YQEKef9K/YiKssWxkZ5ds8SjwddpUfrPx5QjW5bMC4B8i8r974Nqjzo2Wd5s1ykabs6BL5hSwKF5
t9VcTEhr5/qEANTTxjHJUAU0DQ3A9iPgFkeqK338d2w1torw9wFlwgwXf2wXYThTnaLHBLinl6B/
cvBVEPRIpVETk2RmR66acnKpx89DyhiY0Ecdt7pBq+m4gPgK24dBXrc77i7Yw9d74j0MvbnlF5tu
HkuFOTZOEwW8djcTaimzdpApSHyvSxpi1pMDm8kc71Hcov5AM8u7KzcITPPJ7eO3XVpv2faKNd8R
qnLsQ+TfNJfWuORaiOyw5AF+cWTg/SwOrNU8Xpp6/E8xY9WS7IM8HvxZ2sYMOIRSaE1IUf6q1G6u
3wb6Umj40hYycdkUjQcSIAepbGDrFtKqZBvokgyBXFfP9O0S61MEKNxT+wkNBcTpoxZGkwZ5HGKt
qsMnpiJQSNCHI6OWXm/L0cZH6t4G1SwwvFbtQVmqrQ6s3xxFQ9ItjjBqyfO8uKubHTBPRYTDhpau
3iNYYYC8x7jl61qpiPaSo3nGH1B9DJvnauUWB/W5udxNs4nKQ8DHtnlzUkkNC4+oqKxKUiB9WNi2
2EIgAvK0t8AuejpCG/HkxKinC5YpaF2aDUiDPKrq87BArRy0WPKHGv0uO0UOKeZnnsZR0zMayQDE
IRYzYa3sdsvsmYZRrh1ki80A5c8UDSaQ6NJnQnteBKR955AipYJt4TnQc4T6ev8zfmMJKuCZ5thp
jhX3Hwg+xC8EOSguTL1ZSp/uuvdvcOULG2Q320X6PBoNqGWZaW4Xp20s7uTFGtdyNkwO+/X2c2xV
jNDlx4Xis04w/03MoXA/QUf/Z35CeMiZegeaIRIA5F0RE2aK+z4lw85H1OuLeXnohzqDCZE2jkX+
7lYGTAl4bvaN+2MIoEct6Cn+z/AliuazUOcaNP2i+Gusf3UJvCwH1ELwpuxKhR+qZn+HvwfMRcnC
f4YWmixbYwYvV2Py7FYHXAj6ui6OieNfNX/rAjg3K+9HYgSdtNCltkhWdwYhKBbQaryT7HdbpcFZ
z6dhW1OHWcFKJ9k6PHiD88xKlFsyynw6Xk90cndj3rKRYYqlU+mRIWD5raTgX+HQJJ6Y/KKjs14M
1kkrdmk7Y0USY8aFcNCJC8aIWQx9I9b6OEZP6e+dqGeHufcEBGY/5dgZBXw8lL07ScmtxOhuKR8y
AtIo34YUpYD7YgqA3pU9G+x6Ekq4dYtPiH0mG00ZoL9tqzrygvNawpy41KYAkCWMSyUL/eGe/tdZ
Vd6YuFHzQfl/Z5ph1uS3hzSv0ZAdkSxTuTsnQr+8sWz/mIiTuTqzFDudtB64LXUoIOZaDE8s+TVl
BZiTifUCsuItDBZMC1CsuPF2PLSaB5hL4gJno4w6srEjklVOmwbvLZKyVHHuM9vSxc5ov9z47+86
MU2KuiXNFaLhvuO4rwhJsLUtOD06CGGSEyETS6BMNyPZkLhGhtmXmdrAHYIHVXzH7w+pEKTvBNX3
47YFL34fbiPne/pD4a9rsIe6dkYG/ARRbcWzNRoCH506M/TWzXKHmqUMWT9a2u2mrG5KRcHbfEqJ
gsxMesHeaWU6FiQ6V2r2PsfR1Yt+NkS6srWNe6FUK3BsdLSM5oVoo58lVOe+Q4nHz2iS2QFK/2FY
lWEdLPUGmOW59Ccp+Y+0ioCZBFNb0HNM00dhWO9QinMbRDMdIhbt/FaxYqziu/IbbAMxc61V1jVf
niyUxV8wfqxLGfRtImP9xUu+OEwP7uqbb0QblN9zk0h0VU3N2AajiI5hwTap3Fp6qGydSfdQq3Uk
g/PWI5xPuO/J/up4l6UD6cFTMLx63hESukdPcffE/rq3B58AaiCxZ52YUojYY+nNBX7jiA//ZU6f
vkzRPRjiRnNnKrqeaLT4dLQWjinelzwCbWcaokTvqO2bqhggEf1GuuphtJznjDtp3T9etlvA7me8
STi+YStD1QEgHDoxSscqMnrSBw9+UmMFWZjIgQ4hWsp2DdMZyJugYubaM4eLmJQBGEZY9LXkFcYV
YisXj4upEWOoQHPsUt6oemzIAHlNnZ5w/AS9fp4PQg9vZ7ackcrxXj9m7/8exXsLOp/FdNHpjdrE
5mr5vsLpNq3QEuLVreLbZVWSJsexKB9KbrOPWmOXP0y8MviqIE2ssEmk/HxK9WI1Uy39hmnx0LE4
VmDKopImUICBdWvKtyKgVQcnUQXNZ0fku8tjT77gFyCKFGKmM98wKFB49qMOZGzwHzq+N+ovTE7H
SijuJog8Tdcr9d/eLE8qc2+DTgVHfxeCTvS6KILSuKx0z4I7dBV6NaPaEHCKilwq/1ZGxvzXOSjZ
+lT7YRgE0oXGQkEqVTENTPMlUstOzYAepthHS6mbVlFR9i5Yl/CRyUwbGHOa79KY71L3Esscpsb+
19O/uhsLG084OdCw95liElvqMnYTgc0MSYiKJMnIdHEVgZB6c6vYmXiTHoRAggUn5hkZWdfaSYOi
YyXc13BpM0cZCVsZZpniJWqyfnGY8YCgerfOI9SQlN1022hYH19PtIVpwGxEYFdYbAFcN7aKCqpL
ZT63XoxjAgwNb+YJvSMDCu23S9OVx1NOkKKsRC2F3pxPtlCdbC7LtyfviAC1/1Z5UHlf7o4sGQTJ
FJnZrHLQpXaoEsbDdv8JNoHXtXPzGTD/WjtreXTcAcjA35Rq2uxDms1T6iMAbXpPygv4UeDgzEYm
fsrg4JDCXKk1KSVAPvpbSMyTHY0LcWOqxvEou6I6mWFXFnWBejraUTlbQJCJt+fAr1g+hUV8gUVS
qG0QVYejwPv/YsHoq8KuzxXFYxGFiBUtGzRxPn7cGP3Y2A1veWDhVpUqy7XRNSyQ4PYtYlfg8US9
cZ9rNDtIjK8d6viB9O4phDfIOovsLrsRepDiN8GI0SKCJrJ2rS4CrkzBMqyuy8iU4eakKgVe2bM+
APtJVaessLC/6HWVT5QmyPV3ywcgnTIUX/e0MBi9CaT2VWs1PymoqNd+V1DAHnAoZuaZBC+OlzEh
fAJLY3NHZDyI+ynCIoVuvioqnOeg8Dh8g+qnOjVWyi7npRF8MR1sPe2xjOQAwp2hE0Q4+jcRWsng
7iH6gMLRtOjHcQTYiGftZTZ0sgg0gcYk6qMLTKl/1PYAKq4b1TM1qs6kUyLuTClzrwNPG7Xd+/66
gVDIUH36ZPLtGevX64dByFcf0r1Ke68Xazzk8W7Nj5Kp6J+P6wHXPGnmGsHSmI/tlGb7j+CfytGz
C/I4Q3Jv+ht5b/X3z709v+HZJ9fumcSAKP1t8ElzhoZjMQpbqSfSoL4I5abgJDNUfEMYTmolq96R
OWHN2Ah7cMH1rkU6dDIJA7TDDYglmgq5BM+kCuCJwgCLh7EsdzarZoV3bYiXYgJBaW/sBkSYzika
IXC88q1eqWwamjE+k2suN/aS8IrHGEXcz5cb5ynOzx3nmnYVOvGg9OwFMHUQsEmGi1IJmuVtXlKi
mpeIAjwxqz7IYHPFSP4pHrrNhxEZCz+UVBxqx7AaGx2AMsKypXs0imU11mpQlb9k43vgP2FVcdXt
42igF8eg7A7aa4uSYWUCdH1LlTQhFy4F4UZc+PEQbqwmcynOkDHYGHP2x/yIaoujxJUZOmfdSKPH
OVBO/jC4QD+t4EY5KIo+6GcUvIUc79WmF0CrEvy5DIU0smNeJ+G7+9XGAtjJuN25cHvSkyybHh8M
TgZIkyPxtamEdayocSCvQmZv6cDUelRZo5rFJ83LohYVxZPwhBV7vqijVdzEqLul36jEI8ZZ2IQJ
5b+MdRQ7DT5iMlNQ6cWFPMxdj8kz7lBfnhOZy3p3/ZFd4mwA6DLghUXV2DH9e2vqZVo6WICPEB2l
ZqEtPmGj435UiMdp3JXiBolcnFSEPKtifeXyHybrX6AJUq3StrqcDVwRpOlfhXGO0YgdNMCZNa8D
fXckDsK7LT1jrr7urBfXk+EJ372RKxal1cQ8No/K5ftn3rI0fGlAEsLwpwhoDRK7f3KmAIqtuy7D
DnV5w3oqviDFUIzSnQ/NObL5Yw8EEvZEBez6vdAYYMntfMtJDsADeVINwfPmyLSqFvTOYF7f7lD+
+ZWBXhiqAwifbhBRHGaKHFDbX2XVfcyBggJy0WQJz7jw4eDcUTfzj17YpaSs7nODCCkuiWBKRYaL
6bZfMQfARz4RRyMW1DV8PSa+CmkHLS83p6+Z7T7whJX5rAToHMhMXF+92v1qR6aaFP62j6nA5M0R
4R+csu2pyklKbkFNlsJNhaflHoJarT+Ae5/R+05Ym4loxpH+xVB/RNapZG5WUzCYbBWW2IDMp6Qp
NeozO7hJMtxBf6vNerVkJI5nXn68KNh7HaPMyzgFPPRuj9UISYQ95k8Abm1ddiAIDprwTzNHNyWt
b7cJwJt9IZZAjW6JnhPIlp/xRgKp5T1+rgmPQsFJPDtsdQJWHuXumMTgBWF2yzD57sXA2WxugTx1
TqvYY3dx1YQnCqPKSLZ2T9a0XSUwfUhKEA8viFjfNkS03TYrgrOkcriVzHO1IOcg0Whof1+vYnHV
8kC6vaSVWkEGQwqZpa/yC1el854WO2gxSM2NmxLkEHmPHAKK5/U9/RIqWidOXgoxahG+7aEbnchm
HDXFy1QLEAa1jKGPGyWj0tvnfneV08+8lTSYri6snTu3wG/kx8YLI3AVd06Tc7euAGgJYvvNzLJ0
KjhobH0XnkxXgjbHt/zLEMd2S7SATQVRUzXjlDj6JqyySVtkR880q73pL4C8pbtiTq5T4Nf7x4ef
5oR+rrMSpttYdK6sRfozJTs84hnceT8e2F1chE8VCLEjxwdYaO4+VdiM7TiCe0OZtNjkvTRv+k9G
76tkKTq7c+jFtBC5rl1Hi4YQ3+MyG4B3kV+oWIRjvpJp0hpEcqhTWl1zaxOm6egKhdi+wmiISpPM
rWBUJw6k1m8k4SuNuOj346Q/OcU6b3qJ4eeO1OnpBU1wn4gsKi0WZQ0Rly6SS7UxbWbIuFZUomaj
oOr9juOPIiq9tiKeMHFpXr9+sia8D9sYfUdbfWC8sYb/ICXGxPdcIPuF6PI8qCqpOEoom/yDMFj7
f8rgE50PDNfvNUzLOwBbDxg4KhucqG0Kg0ZqtAXsf6El+pjh8Jm8xjbXDLfWlDMLeHzJ4fpDwznL
/yKqUv0WCZ8jQY/vZsFsm5qKrR2srZCYjXSmu6H8AyNxZ38EJaGFpD2f/I0jl5EIvkuVbzcZ7kTE
AjcbhPPkL9ujjMgPeViCmfdJOeOGUY67C4bsL6+s17OFhD+UYrn2C2S2Zn4XuQH8x4xi3czWrxSe
b5lpyicBEbsTshqyX1tVc774n9GdQjijLxIqGpfYIO2cVK3fa2bLymqz109EkoA7MyE8Movx7rDz
d1qK0ZmTOoSrd3nbysPVtrZVEB0EwoK50i5FEBQNkmQ/gzEvwCIM0wsoMC6KGRdXvAAOwyM6fmRp
AJgt+CZHUqHPr/mVONRGsLrLZN8x+T0ugCntsVU31tQEWPJLOMFHiHMATixdq53SLff2zBDQO2kO
nBauJzUevSHEYZd2q9pHSPbQ0jMRLosiBtaf7602J3SGzbtUv/W8/selj6nNIbQHFt0P3u4OO+MJ
hzoItFE/X61PYbHgy+9Ez8ELBcWrD0WhYC5KR3WrOtXmYxPxTy6LY/st71kB1udQ64NkfA3wZx7X
TMSamY0gze3bkdiNudwuxdpFA5SCVN4sL1SC0GQpeyW7W9anO1xBpqhpDkuFhFfqicn890Tn5P+Y
NM9mTgkOdm/DpugSQqTsqOb5fo9oeVXj5mmR2g79fvcSydhU4U4Jv6plwcN+118lGR1XW2L04PA1
Bnv340BjeMhjjHFoB+1C/haUghUAFSRN8tFx6C1dK6KoJfxuDinm84nhyqgwX7JSKgB7U1pPRF/W
ATEMmQqSGPC8kNaY3KAJe99tyckFQamKbXIdBfzlSJNw/w0KoUbpIi7p/hCXZTYKqihhjs5D1EJl
3owWS/hf3o6Yij4lOuAT8DhNmoxkXfFi5LrLA0uOdqxhkg1lBKLzcWtBOTmP3nS2fgfB8Ffo7mZx
cE5QckB9qIPAEk85G97A4oBgSr0GhpzT5n3ya9eRyAkdwpZ8+2Ah2qjt4Bsn67COaF37pwwDWFkk
Tx77EblK4DY0LtEKB3a8GbotQOFaRzuD+yEGcmeldGEmST0y3FUPwgxDJLYUsNg5qfpzKxeDYFny
Iqj89EYkcRa1xvGhwgaduSzUkZeGKfRyDg4pVz5s/yIcCf60I0Te4OtIQcviKMrhndecAqAQ63C5
HJ6raE/MnSnWbQ+KOvJX2+AsQU2JDWi0UEkCt2Z4XfFFkhLJnuDV4dMw5/b1Rauk6ynqCQz04cIF
hhJUlEGgWggnCwgPUXknETg012gmfolan8RIvkXU8h5yOnhgNCbXCVEHJ89WgmAbR3t2sNQDjQMa
U2w/RYAg1SzXCNbEXNqvRdAR8DUfGcnbn+CH02Omx5/6JDMYiXSBt+HaDBO9ZfQpFsR6yX2TGz8D
0jworGowtq7li9hp2GFqxK36McTI6kmHVI39Nph7Bwyw6vbTiNWjTNs5W/mr2hYzu3opac0bIHx9
kC9Vj5Q+xGMBWIw8G/69W5dx05pJhueqSENeU8S/riaJZP9zM1B7uZnfvEcs3wQOU8DaVzukFJE7
Kg9yRSA919d8mvzssLqp2G8wtEd17z5Gu/E92fX+d7wYz6CtNMMj7ym1qB93K6EG3SRg+qUk6CcW
V4Nn7JTsObIrm1ub1pKoKg0752A3zBEpSId1HNnjJxvOZ2yDmsaNXjpGxkPHlPu868Sia9qx55ZO
ArrNDTLFTbuibyKqSnprJ7QbVwnnI0P/GdkId4rhR8bT4w/Y4//D9SJICAnDURmy/kTux/6VXFkZ
minPwS2GDscztq/vVc7RKRaG6zNOylfvhyUdtj5JaCCEqJ8dXk+RKKjHeQzU553ShW7TwcmusRGl
bIIfbqT6APFfF+tbMoET5A1mjPqnX9+ml+hy22nUQqRwWvhiLz7geH9gxRMYD5bcI7xavajnhkJO
y089kOHFCiMieyoYoAMFqbaDdkf2RWiwoKUdSjqxkC/nwi4PD711ZpQ9KlPJSyEPSU2TJtrs5vn8
+cj8a1qmMqUTC66lQCk8CCGyaCt93u6WjvBXHjs9gDBaoWLKAlIETf6fMizh5b8Q4W0p7XDA1Yxr
1p4YRwggoAXopj2DtHIydc5C3SdlTqIkY1vXVwqk/qxvyFRwnJiErV46eLbww8NtutoNFRBbZWL6
sUPg9J+SoqXzphQs78XUon+3uWm8yktDpGIuy9f5+qH8SFYJXXHGr+J4bbK4aIKkCu7GKj2IqUJH
htwG3QN+R6/s93LxSGzkBIu0RFLjcTN9Vxxd2XkVSn9ChWzfbK9eeBBQpZcpuGfEUaIrKwyyHXeH
hLFEMIdBK5B3MC+Rb1e0QC3xRflmqhQi+6tBu97F2eSGbgrgQDPK6NLHRaXjhqEEIY06WYO5MJhe
MWcPt1hp4rqYT2gbJVpS/nB0DqU27Wz6SljIu9lzYh/ZzfxNcoxj7qKGSGO05s/of7MFJn7Dn8WR
Ur34zTLnKjZHSfxdNmp6jZ2tSJtEDC3IqUOHKlOCsINZCCSO64lRH6TuJ/+IU5sgDX/4fMizLlEG
q1I/LjITABj1CxmKq6UZqnPLLu8TfeTs2WehdwQLutXwtKpcXDu45N7dgAVN9okawx7LZZNoeO6j
W9sWjBjTywMzOSKOFsHR+HMz8zvk66Ih3GMyo+bPuyH2UTH1uAQDs9Bw0SlT+OW4N+bpR1vjsjJ6
nwtv+oIYtmibAV9ax5enGLD3eN9+EIToJeG6HkOIrlt267UPYp1BGkZDf2ImGU+05HqyhPsMnZN6
7YULUjbEY8kNu44PEGqKttMG1zJV23d3BjB7/w+gt2ijiEbIRwNOyOvuaVyV0xAbqjZbwJRcJ46P
MS8Q8wDg1maoFm1yn1EbNIB8eWzYXyW3EJSTS8JiVHSCZHEcXvPaYQgExugy/W7uoIgxAf1eMpDs
8ym8N3oHVtK1bHXubK/BI+EGHnWHHtkxkQOYvuz0lJqNeONDA2flmElKoZisWRRoFgf7cJy1+Tp/
TnsUtuvFF52dNpVEjPdi3tYG701roXKzY+rs19la3JaOtcRK/4QkFU3px1lC8/qOdu95X0PjEQK6
yuN7uAqRpC3/b7Pv7BH0u0sscaxkRklLtjnOeZScM9nxn218598uamYTe/uzZX5iPnBEE5bh54hl
9aaCkiDURnOiNjWhWDv9YxOfp1H414gUpr9Sj8NPGWXUctJbQhFWk9odQT+ylMGBIpYPaO77sS96
WqrqiXt8Y/7dgGtwuUtPRwuNQcpfU2jB0cTeeaDB+OvHspWH2kz3j3bHh8rbIIwOrwUSKEwLwi6k
ihdY6TSbbWEz01mjIXh5eDNs2UtGVraQcB7vX4cqS1L4t/jwhmWR1KrK4pofX9tE8PQTcUdpBMK4
+sb9FMemMWKIWVUbG0lfT8IRzPQ+Ry5dNku2uuUArJVRHDEEc5yLd0KzSXulNNbPbr/6J9vbeDWp
5ExZ/QI7ZcwWDoT/6Oj5Ue/pXdDTtg9VBHkd1NKvXTStwB14DJ8nTftRaswnONSssjO8y1e4Q8tt
6f17OG6jLLYpHVs02Xm4pc14sZWgzXaUZ6Kb1gAmSQZtmjvVnWfYj0T0slvbZCdP+4/F44ocLrMG
SmYHANx/vhDL0DdA1V+xXSCRJ8wc7ieWPdoL+BO2P2AZUz6f5U++PxS7WJty7PvTYUpJyV1n6OPq
QwxlG2fuRnzC+rx4vV1CXB1/Tjw4I9zL4w4KAnoyRSHjvemFBYLWaJt9/9flynJ5IsHy/IpDVUoR
UsLK7srviAX5Vce7lzduL0isRGNv6jlUkXygrglAhjixM+VpoNT0JFYRxFPaUrN7ZJtzh/mnR/4a
sbwwZSXHqJiSIYoGfbrSEoaLKI2vMmOjDvRf7eCT+ieantogp/hNU3T7uXb35KF9v3rcSqEtx0/L
J2dkB0OzQR1Ipk8TGjjjH0QhDE1o+vjWBdNRGwxJGChMGTZrpaPPmmnjruRaclnKUJpFkct68hmH
Pb8UIHGV4paS1PBKgVztJ0A1KOxltmwpDdiWPOLgJ2hyP+0dxdEjFuz4tm91+hzZ4GQFajofkuZV
a1h0sh0dTjbTT+N14BLzxxZN5PP4H/d5pOi1WLHdPolosF/XI5e0oCL3XP/l3UCi9OIJJBkiNf1Y
wg8V7nyDQVXtGOlnDUiHbTMbZ/fI50qrD8HZ3Ukx1S0vz9cEWPkZCX6QyzEv41SpBhRkizvmHtxx
HnWBHbniOovnQvV+s30RYinFIOe8BgA1oqVTT3pMjyK46dHw2Qn49xSkDWB4rKF+Cq7pf3rAV095
9piHcKo2HHxMlG73hi8+fZnq4lIWcOdpM4IzFqpJdWLXcmOBNZmsO5cZ8lFCO52I+Ez9nMua+xAb
vMuyQajQXJH2QCX56bEp3y18/j2LyedwpGaV5olfDJ7eyRT32NzwflYBZhiaqeZpxCQasEpDw87E
76Lrt0vzrowsaVJm1JJB6TQr1XoRUh2qvbqZlayPeSG0Fy/iU0i9WD2rsWLMGDhD6cZkCvEeY9f8
lo/l/gqaNzJMWkoatuU283AXpDXoSwAA8AQbV/VhqZB3TnJ2eGunrH9Ag/qZaND5oLja/74vx28C
Ar7aG5VXhMjgc5p8QtQR2v51IRkPcok7sISr4TUPCzrhEHBnbvZQHavYCWKu+Y+s2UOMGJY72sza
eig/KPsqkV9HFc3BNIYhfQ1nOsopVRmwbNjSYqSGIY1iisBvMEhFp+6uNG7TtN6nZNYWEeQzfE58
+PLVkXNQOBGCmXc/ZoTqjAi7vrlX+PNODp5fyA0dMyRWMtB+V5nASMPskSYG7unUibM6z7kMl2a7
uS6MizJu2yXpCfVH48Q/t3Ncmxor0NPVoYUTK/eH6eNPXIEQ+12AfC/A9GezVYDrzJ/vfA8vhDrp
8st5ObWR99qlDgbBfxXYzs5xvC9ROyg+Qh7ScG0wxGdB1IXZq41YA425noc4uscIuQ5zVBIHNc2s
X5lKrrJ38RRSH95cP2qYOnwWoZcva/eMhkcmzHVAQKMVQ1yqnGUrjpPY3vhlQLRVCQEpcrQjbjaO
nX9A7t9RZ4nBUGL0lUzbJLDdZm98IwKdj/70ZdsYWPwDf3KbYTj6QeA5U9zFr0UTHpCj7JGjojo1
cyFPGVcuXk0nSpinDAY2waBCRGMbNw0NCN4gNIIXengI94COBL6eIfjbwYMDkYK9TPH1m8155E5W
EokDZn92uimMeGw+vOrwCZheork3SoNBuLxYccEZm3SRdM8PPGLkULAomzjhm7lgfV/zv6/WDdyx
cOhJLHOqhEaHRB5HHhw/zDe6lrf4blB4XHY4EwD08BHGeirYERvABPySV/u607J1P+nn36Ed+Zbf
vYq2AjD1eY6UDEVn/xcbOt5MX05A43Tt1nEba+nzLo7x7PWP1Ht97a4umdgxqP0Z2wJIxKJcr11m
cW+fgcX/y17t/hp+Bgve1qE830uPAQa1stTh+zkZV18MtTzjhIRBd7ZYOxEU3bnuCOQbbCSPMvrL
/ycZoqGC72+CjSS4z4Tsf7mpsW4K/L1z9ab0RZKahN9zx0nFzAFw7qOn5Ly6zkQ7alhIXA0w0hJo
k8BZgdNrLvgDUPReIRKMVBV/4/0sKw8WQGSfruKIAf/zHJC0jfKBBySUU0lKpBSycLI4+3ITFd2f
vWQK7eB3i62giYZszCxSEC46LPJgzoEOLx33Syy6dsVvm1eK92NlYL7hntW9WX1ZF/fL18YvUPC/
F5C4yfmkpqhCr7ebD4oOHDowyB3WZSInDDoHdWYrr4RpD5xnaoLLociDYbQen2GD081Jw1UBqxn5
5pEpRco+Y6EE7FyQmV9k/kZgnfJTKvqoCeICpAMttSqRpfFiyVbHm+/7fX07CUXmGKlnev5a7EBl
yq6fRJs7Qj6iY2DkPqKjP2YSE2+8/YUoX43CVqqhkJIpQEXd+bi32tX7Jfr31nhGsmpeReTJoxj8
AmPnhxqH/Z49tuleCZhj6yH4xTlyxMwIC1r2LJ7VMjzZtniOetzp07IsC+vPsYlWmYcrJ1Y4npBN
eLLu41x3iX83Z3PMgFg8S0AKnv5W9V5fGtHabZf1+XVXSb5pAWJZp3Y1x9hv3GYVJID3wZ0qLfNv
r8ObLo3UejlZ+wAhQTPM7j3gj+GnhXuz5BbGIcJl5VK+UeYzDK1yLGmVAj/i7qcBrJ/YQqADceHK
TzhGT7ZDTva53ZDbL6H7pV0X0X3VhY+od+ANWFv4uxwZVKXFGeae6hcVmTJNblD0kq1iUyL+hfN7
8puhJCHnHUkOrbLJzRjgUrI73hcMDtu4gncK+iyCJuxMeg0KuoJwnObUZSqMLoyzZtyX40KjT5vv
3zDQozhrUXNcKamt5vQuBGzNy8IwxWfRoSTd5VZ064VVJzPkp3GcWD37Z0KNmAjTRM9PlUPZohWF
6My8wRqnDdI1vOtMPw+Ckkka9uwZPhyy+fYyP+ps+ThbSo+vY43+2kjikBX8XueJqMKlm1XDb+we
v4abs8s0cW9XP1K+K8vZlBC6mUDPIqd85B2TnEnNR4a+8YddnPGjRrEQorHHIfXjR8t0iPin0hol
y4qL4aVSjxE0fAaT3A1JTGEB2rcE30x6X2ue00egzRZ1PMplgFGvJXCnn7QCBeKWPjL7q++KKr03
ErYYdXOmvNxWsTz5mDRLgm1lFoFHf8Hvkj8e1oewwIyJWGOpxCVQT2KnE4DiO9TKp0k7cBsa6Eft
uolsn57+BR3Ymns0Dhv9drCOYLzcNfMRE/bE8mEfs9KKz+s5BS5yj4111djUDigeKtyGVndFMv79
quGSw5JK7SWLNbEu+ecUzQEBwywb6amvhdMFFTlO74NkrcKvu6DVtzZg4NFY8KkA/Sn0B+VPdSgY
BDIeUVqoqQ3IPBAjhSRWIBvcOHDpvOVYAjmB44Zk9B6UcOdFxMugsHF535tmLbXxsb99woFdcbIb
3dh2GqGrN+AxEfJcIpTi1409qk0u9WPEXe0eXQeiQI/lXKV0IifJMfxWMJcPiSQMa6v8R+F6MViD
7nFmcKcupKQ/hQ6G8X9eiLglQRCEwr05IFs/Maou8qG3eMbA+7IEpDC3BdabbWOOZez4SEG51oen
29LN5LeiNRR/GT3MYHBVqUtOsXxSnq4lWDcxxnVGKZORSCvtEfPuQEbSLDhBO47HZdYLtz+LaAgp
TzAhGMz6Jw8KJiY1OkRvJ69TwskZfC//vhcrXcDvawGMsaHFgO693qUVwldShsw4bhrZJk5WdXsS
sxrzaER0sDxxyCg+p+/4518ZedMucQa3VMrtbWvstmCPmp6A7XoHYlWq7YBtqEHwUUPEJ81K8w3E
xvVDfJ/JGPK0KRFkZc+1VpBg4GkdN6bb4UkUe40gF8v117k7+88yBV3ELszYEvlkbMtcGoiYOiB4
o86dnOqFNTC95nW6rHB07qZDVk+3/0evIcJNGEoVOi7rvnGnX5EdIsHq6WAKVOmxB1W0XFbxRCG8
jskDKIVRLIFFlul9tK6en6OrRBCI74OPweKbhQcv0uMnjtnU2S44BGwHz3q4vQsEYqzJrdOqaIMe
EF/CEtK7UgJbnwkViw6TWc7fw4Ybxw+z1kKvx5CwD/MpXv5+yEbczUpNooqzv1KV0iv9SBwGalBb
swjjlD//fyqAO/3+RlUeSErjR86R7eF1sjsyYd26sDYtrg/4NbH2rNkbSwAKPLT4k2InyPSqEem5
c198dpjO3bsZfYjvM6wxj6maVgPO/x/iEcqltGlXgekikm8kaTkm9sCnJhMhmZD3SXMcfgKze8S7
BuWA76jw1qt8khltowBh9PGnXQHfjklxwduGaqw21u2dIscmJJuzPRYBujyuEp9clVEjJun6c/yL
c7tuh2TPQK8ScFzuo/AGRPZUeoNqXmn44bW3ADn5oD9JaPsBP98nLRSEPVljueMgWZaBck7CQKtA
QrG0F0W/C98YjkPjMvCn9aYzCEkRAr2kh3WKXAtXClF1CSbTUk+69h8Z262tNn6WL8N66vWQ22YW
KxbJbBDBXzqwFtYbFzBlmeO81O6jAf6CA0RT4gwoViSddpsF1H9anYWrtHi+yqIPdw/lTd8cSgF4
Jr85EYZP9Lqr3B1x/bJ5g9Un9m84aVq2eyrTfZYPia9fc0IfcE3thijcqLI/G3x5mW8bAUzP0oL/
BULl/FiP/NbMGx14gi0trhRJFsSk3dP6l2a2KIpX7m4j41MEw9JVoAP/5jn53fm5lPzb1g+3Nfh/
5GdyclFxh0yzRL7WD9kXm7IeG1JrCGwyjz8un0YFg+8nQssUB0HtLbb50ju3hmDlk0B86wckXP1h
KzGgVB3u1hxoD4GM0/bj1tfDwD51CYnLkCD+GEFgcK2J3T/c+21ovlLAzPuG5aw1b5OVblEfzrJh
8CcEPiQzugJujkK8ggJfKfnZMI92fyszoZPVeSnlQQrNckm5xpSHrUNd54OJ6dKVwXeqpBLsykSR
/WsOcHaHHrDnhOePwKRMeyHuCkLv1DWTrL5roTx5dAw5icrQCbTg1ns4drIQt+3MKiX1P5xCnYoa
Bc2qeqBMmKfmmVDsOvElyNSoiCigOL6s/Wr+veuz2jC3mpG3gt1u+WNd83uMBRdj6RMVMrs6yrSC
7UKELLxlW3jM1GHdc8tLVzE3/aw3dApHj1WN0mQg0j7aLzO/iFrU3jQgh2T1iPIUcMHTEAUYedOF
D6FszwMMldQ61Y/uvZRvUFW3SUTux2U7xL0gy1LdGZ95MAqOXz31/lJRSxrNV7Wz/i7SZVb7cfNa
7qH54gf8LwZmewLSV4Udcxe+lGKjohtRZzqlr0MnNY4qVdP4agmSvdlV0UJzJHLA1z6fw6UoRpet
I0egGxY6P8vx+O89KI+9XynbJnX+aMAYcOLHmss4ec70jd/0/Ck12AX37oOy2040e0hVSyTVOsdj
sdFzU+abxF2fbd9OmovUVJjnynBJ7dS5fop1EROmRBbx5zzIXSZ1vKNb/zTxk58rZXSvq6/GQ0qB
l+hJK5uO87RNkTQcoENzTygDXUetnkzi8f2Sh72FqlIE7a2AC/2C9mL/de0PmDBFth3WTavXsIEx
fYSBHUAuzKzrEU3BPVGPYwpPyOXQhsaihOMRhXRUE59j3P76vSq5idY2tzdqyVqt72ao7tJPX1oU
I6WbNn8nrPlzUlSbQwQwsyZX3NM2qAVZffQDhU8urccJV0a1RDrfat2l0NwOe3ONFW2mTcI6LnWl
hP/7r332msOXtKFeq9i7c3i1LiDzuLdmkB7jv1a5F00Z3bpgqPQHcEqRIdBLesmO6N7E/5Ly9uwP
iornPMfcNWKJKXoPrJmfGo4hPEx3ovofKFzv3vALIFBu/vuvHHkx4FDi1Fzmiy4BTdpbOakuXkMG
IZU+6a69n2b/hjPAPwnQt3ZpW5q7/wPFzve+0J0Gjfq9EmDQMfn4DCO+iMTYNOZN2QYU0l+h36MT
6dozLhjLd3G+2dj5p8nqKG/GHjIo7dUgEtEZjMEedvegfi/3X1+fxcN5VgYlKH+5jD4+SSzQSNJh
QBeRcB/VLJPPyj5OQGo1SDYLNarqfaAuQ97yEiEyU2jcTFu89/jggpJfYf1TSk3nHNCaDa2cKuOe
P0PRCGl5yq7/vX++BkaoecnL16uQaYkCyhUXGCV1vT6Q/puM3AEiO90OodWLUK4M+5/buopR+bDN
Gyz/beuabMmJeeY6C3d7B0P/mLGes3xnK+XOF4QCKNBikazHB8Z23MUIKf05NtOdN9DniBdDZc6H
SqcSYMsHT1NOTE7KH+TweVdCuvIDTKm6id1eqLowUy0jILLEJ9VBVsZ6fSPooS0sF+wiur2etrQw
uYzAQHn6HLBHPMcd5xv59/TAGo6CBZ35ZmBBedaK50kDy4w7jb/HLXD2dYEGoXwclXqyzb8EHqiW
bA/rH5m920MRXKtUbkEC+NnFB/2zGhz3xfOwgPAIp4KyJrMljMTEXXTy0UwvBSdMA6wiSuPCnYDz
v6lm7+myQYZBNfPgwvybjF8n7q8FzltZhUdHGwYpPgmisfoRfYjQt7HR6z+miwoniEwslq5/qjwx
R7VTygdsDXDDFCemNJYRW0BDRQN67DfYC7idC2LoowggqFQ43j16uTMcEfv943uPkPqBVyH3i+Po
76tZyOVMRlYMw7POb7cb8FgloGSQckWUkoHEgZPZE1Zpq1u0YzKb5V1g2PGrH1PQxPV3VV5ag+2b
gm2F9eY4rpFcJk5nCX0zev90yTL/ox8sgkrF4MobPB+mFx4Aa/aWONkl8S1q/uqv01bOOUQSt8+/
mySsRXlR6GkMVQRc1HB0wvFRShIV5h2Y6woPbgr8uvq+MlvwwvnDcUoltC5kNBr0yaAjxGKGbwr1
AUq9he8qDXkuGNWQy9BdaEcVF5GAWaE0Rgw0rmSMtwWAKH7cI6VzQ1sY6MMSXycDP2+mC/MSmW8s
xVrB/sm7k5/I1vTpX/J9uFCc8mjdokJ24sC+c6tTHAW4gp/8pb8a0w/1QR1i/P5UOzZBj3lN4YFv
AvBmh0XvD04z+a3jAVXKS9Zm5K+p/Jixne0SgfixyXa3nl8GaY8eIoTDOJ3hXei36XbrMVqcb3/H
aTBgn0jZjyB2d8jd424OK40gu3hmDUzI3kUqYFQpsx8Xtc5wC82TPAG4Wb4nI3AJaMmMVK4iQwWc
IvajjT9eDLDzKbFGdFfIfOyDXodlpYqZOiEp0PD5uusoy12+JLmKtQUdgF/2rsWjfq5Cw255GVb4
FeY5oVoq7WpMeq6Rx+wXdV34Jb0HAQS6TSOMBKW+VR6hiJTXwS3wvCY5x3RfckdqLEjZ4iOPrUbv
7jXAyDjigh1vJ9r5b7T4V2vCqBg+7xdftklg5e6osB3IZQRo7seg7NbB1Mb+Hq9xeP3DTC7tKjtE
zSn5z1JMx9QX5lJRzK7IAxvKsCaIo2wFQKWCoPze2WhUDbo8BovWnae5DmvhUW3zcjTcUvZ0khEY
vW5PqIzzGYmve8KkwO9hGy9DAohfuZo0QbSclUFWwJ8aQkBMzFSW8Ma6vC1/f++RV4wOm/q4K/Kk
NtCCPdrN58e+S7OUHJSmA6YIjKFEOF3KRB9e6cNWUpjtAgu2BFYiI7Jqh+D+sSxZbu9uk4DUYp5a
lBMAZpQNyjztAfJlkcXFpFWdNQ70V/rwtg1wrKDVx5Z+lZuvafcZnaoRyU4dvHcsUP6VOdoVitIi
rZa67L+J2WYL114L5psrwlvU/HcrS2m6yxUiSzmmP+40Kun6XCcgG71SYGJCkNrxDkmbEswaoQTq
HqmQgZ6MUWYwyNUXrjGZ0oG3RSPesmcmStXYP+6IeTVsQxC7Lxe3Iuxbjst15kJv+BVLVRgxZ9Gs
pjn2yftyaldQzxaRXsaBxJbrD/UxQ2HESjpfTl8e8Y9xpWj/rH0PO2Pk8V5rgDbtEZsAZGp+2iMr
3PThWhOgPq1aSKguVCmK1w6UXogehcZaPnaXleEcRCTEpybmTFQ2HFggBUYuIEVIjkk4R429zmIM
UeSVIgqts9UO95jMjUe6Exrjd2tQ+FXZtqUvVr/6RBBe08Bdht1ZGWX4hg+EYOL9OkYXu5ZzxQxm
dWrzrZc5+jwfLGZxmz7qZ6PrWAVrqjoKrnFb2paXI/oR5yuclmRBqtdA/ktOAIfjrPOwGiK4AT9h
M3nGej3tHILsirA3MvGv6jAXrOU79eYXiIQDLgzwMUs/RK2VJppLi9Xg8FTTIOJoKTRSXVepDMSP
7BkJia9wLDE8WeZSmhfR33XhD7NJ+1wPLVJMR6/Od3gZwcNCXccTU2oaStDVgxHlXGivIgI9YeUM
gLe+0LcIXHYTSAWWjkrewBYFJo/oh61+4zGjpSzIx2B7tDBOspAbRC9/35o3I5/SZn5aZ1Mgan6Z
K+j3NV3qonMJIbS7DjGxfHR2rXQDAA/7zA/eSEqUGjoYitRMxwBC9UWRGa0sr4umOLb4YrOa2QaI
E1MlbHHFRl62kQDzf6p+c6HW5h8EAvsdiz0d9AfFvqDC3YVlfSLU3ojhIfONYBDcJTDoUhlNKZyx
uLSd1nn2j2R+MmohnPpG0U6/lanaPB/9W+yqwp0q3LTyglNPPZVPH5xMNUOw76fsuQbTUTUl2iK2
mF/41z/PPX4jbiETTyVHPaZDMAE9eKTKCnfEGeYE4Xi5VPsmO8mnBLn6V9ttDDsd92W6METrPq80
LnRMV/eh8p1vCqBeQGSWCNE6FbufqBGUGRzNKlfd1cXOIwY8XaZSraiftwxhBVjv2jBkEm0nyvBS
ZzHfETPchiPA1NaF98G4jy3yfZHLhESPwPI9KIyurTYy9018LWBrNwVIO0Y1E0dPkQAUJ46CDqHj
I2zmeClDUGQirSkeHHjWaZygxdyvjtsb3g4Z1BgVlrCWojaO0p2Vqc3G3Rpt/HF+3us4Qm8esYUc
k+/r+fEYYeTUpkZ3dL3Z2obEKuGOcI1g1yABlwrmGgHkyoAmCMBjEXiSEtgpEmEvns+Qryphq8g2
49M06fpVPsNBeyEguGDifDApWBFC2Koio98Pw2ulk50/X4uuXhixfMMQcVCM8I5O5UQW7QrwRQtw
xNrbf82HTcVdEEsFQBQOyW5ENF027YhlWpH0yradAeM9haiOmqG+NRJiSDnIZTjkePlxvYCDJlHA
mzodXd97AgY7tUi7FTaSgdIVeTWfe6byFJOVl7yK2gjVq2Pleqf1QCtIh1R/1JNs+ulhs8nSWzPo
pZeRsjeuTmpFRFeHa00T6NEtSdvC5hV3HUCmbEY+T+6qcju2SQ6OzSi9ICLQwWdAoIQloskTjFm9
eue7sinwkiJOxyhFBebFMistvJkzoBEGz2dlONELc6LHKCWdF7Mv1Kp3VNldisF/X+MoVgoGdyK1
W4XNNZI8etP8yCFHDYU0Gh988Jory1AH0GYVLCuhapIhXib/6Jxd0vIxTAHtt62qWEF1xcbNYTnv
taasF6Vp1a0VK7TsKD4vTIsK6H5pOCevkW2vthb1x/t2YF/JjlFoU8G49NeARGqf8rX2giWdXi8e
s5kTh+cCA3+s/WM24E2OVqYHSX8c/a4dy/H2tmK+LAdHDhkGWJRGM+jdc+D5LHGvUb+tZPeAVKLP
t1jEXvWSmwPaXRHlfv8iCrrJK8AOs+xX+0oStwyiSsjwcezPOxSlx+0s/T48CkYFUQ6iiZrn/Kgh
bY6KDH64tv6dfhJSgoLpuUQgDiElGmVPj4UbiQ5uuw/CGxEVnW1s1Mzalu4kgmRBIHZLzsw6NUTA
AwQuuzoSGaFP6QzmhryCrF5JDh6VGeFaYdi5/+NuZnQB7CvanNdNh+UMks8IyhtNqQYh0GtOqkwt
7LCV3Thwe2bD6aua7CYuYpIbFHmWMZjQcx8IpzrmWnrYXhlGR2dsHVFPOVP5u5MbbVzjTVtfpjmt
jwKhMKhVUNUv06HpWKjX54uMwyR65eveSH9RQiggS4ddkk4uLGQ8P0EmLdwj3fMZvDcAM2dmF2hL
vYr1eXimEjdUVYeNkvVs+0w2am4+F1rV2J6ncuv1iWTFXf1IT2chebxuMX/JW1kyaPzKwe91rix+
I3ronxk8snkPmQtjziOaKxpwk3GUe+m/M4fQiba/q8A+7c73dAIXy/W/Ow65PV69qEchK1tI3+xj
wnPg+D5C08pmpSpjxzN9mP6dO1LpGP0LNg0/zZtK6vLtmSAkebvIJ9gfslBerq26T7fPa9kfy03P
h8g/ShRCN3scVfvpVsUmjGF8uQx/FRHIobXI1Fy2fPANmegMLvCGbbdfDCTeuhM54+DmaUN6+R+K
+oVkbXYI2T/uCRPM2UeOhz1kyGGu+BY/d62ipsWToRBIz/iiQvGLkq/ikc7hVV/ubRAnWLefRqyb
q4hXmDvGUw/dFlwLS4+0+cgONOUbA76lbSTmtWPTgidsOmMnd/68iQFmg4iGcCdTSMyh3nA8V4pq
xBmXeg+QrN3GQYAJ7GWj8v6XNnrwVCyifJuhLIDNu4aS9aF2yg1Bi6Z3Xoxq9789/b1ikOGlR+rp
QvRRm3g/pq2fmqmcA4tO+BjG+OErLj1FYtiPrC/GJdqKf05UvDgSP65QUdhc/z4K/Kj92TF7rSjg
c2zYG61ycW5LgBnjrexXv1+qON0nBxCEHUjATaemU1kIHDwo01ySO4hcABKJhHapJ52oxt0c48+b
q4HsVBHJR8hU3ClnxWDzX8w1Px7HEpHW2vIl2Mg4YDy/NIMOPWkrYoa4IeThdkL5YQVllXyzuO07
NrYQqmkdlJJ/AADLxr3YEXP5rE1tf2UeYBwJgJWx320pwPnmYtOKy494JC81s9IyJ1urbhwLmfvJ
XCeMwVUEY593ojQ9ONvtT+xcoYEgUg63jtCLoq1WWzXTTbkYheAbPRnmXwI1/BOWFyt6/7F2gQ+p
2go2aLU+kgWPnXAzMeR7WhLNQ747MuKG2nQF3EsO5t3X5++H+fh84tjeg58SJ4N+nXVvyvidKOBF
oN5Q0+p9qY9TauDWvCiHR6DJnUGsZNkYR3/j1Tao6ULgZu8sjqPp0jUo/Hz2hlUFzstrid7c3ezG
fwFkmIhrhidv87dlOJ7I10sZrxXDXJr8mGrm0T+qZLgZ6PMHsHn2N3BBny79PPNpr74d8l9pi4la
Zb9dafXjQyDgMmiYZy9oozO+0Hw7CH/rcN15kXhJAWF7TLQHUls/N4hBoFu/P/1HsYKYJs8xHQbV
yoisCOxJxPyxgTVpXPGi2bpEXG/lvTKUarLmpzUnMEdX7ljkamxUVTzH2hH34xELfA+HSchP0lbQ
h7DzoN81PXV1PZHILH5jajavU4B/TwEIb8SyAIwDIg5X4lrb7j1yr7yx6ls1NN4tNj0DIWtOBDbY
HsHSseY1UX7itVCwkKBnlkFd4VsA1Eye5MzW/qTV46zPbGdJnH8Rfa7nFStHRNWDzjsgsu9ytSao
e67+Ice6D57BleCNj9NbG3hO+mhLR3U5TGAYEPpgsNoz+4bCwT0Qf1TSzhVOMcMB2xjau38aPcK+
gNeWd3lZCpTQrnogV5rabx4LvKMraPdSLyl23lunA21YMCQjrKWCCvAlP0Bv09qG9LRDVRjVwS2Z
atRS3xPwQpoR9Bxdw75d74T2sfCwQhK7mIjwxBWlCPzJ8D7JSNCHiz8Sdlunvf4Ht43aqmmJi9n5
QvRQq652GgIxRQNHcg/iif1zy8swV5IvuciN05PDbLgSHfhcyGaezNs068eJ/gufWzblYZ+TaQ7T
LySe5bV65/qUWriPxs35OYyl8kg5FKczbH3StGnt4D3TykS2DTbADl72hbgspJ3AdbYMJAwZINkL
q8XR5tFYFqFp1r6W1EYM5oHp0hCBj5A9ps+SZ8A5DdS3b2HIy9Wdv9gWsKyk56eB2iZI+It1uVQp
1GETwPwM/35f5IM9qceprayBfRZK6wU0uKAQoYjUyKRXY09Pc50szooJNF9fHQSmY5+UW09csJUZ
9m00RPFZOS/f0TOW4No7lYB9rm/ZYUppGe5npYdhWHd4f4dAMRGBxW4BXyVexw0S16L3UwyVTFOz
Vjq3qxNQCFfedxV7lvll/oTDDjCZOqCKiS1a+X+N+RBGWWwoBcxmM7aqua6JY6vIma0wp7y7cssD
2pkKW5MEcayyyu2NNOefMfP5YBSByqRqRrvIOQH9aj2+OoSFAKM+Pspbn10C4TrqAI5L6Q9RKmVz
CozzjmAL6/91xA5H9kzeDlzmTvH98UQxCP1+mdckMURx55rFWNwlaysY+5YdlDqlapuTJKXrhnG3
kMrzBR3cJFbnHnrTJudXKn2+OpA8OpikrzNRXfHG+la09tkESxtQrIw4CxUD6eIJOWpgWn9qO5E4
iTcg0mnpOQPH/47V5IK9dUg7w3WHLCG3n/5S9U4u8xL5ZpXU12+VmzPjC4Ys1wV7uX4nfCac4DGn
ox8FFtQPv26OLMMtyvRkLcdKTe53l+sQD1ckdjctto+L6EjmPcvc+pWL1w+gxqQJ1oizyI1i/Jj2
XBvZqLGcF4TcvX1SOWfs/sAUUl7WmXPvBfBEoHXu0XUrfcufhQJ8Cw6PJ+Rg+/KkQ6W66Q5D7YVg
BktB1M5+xwM1djrH9A2M4hKhl5eve+XR1dJe+TLCmxuGgP9Begdr7QfLmodkQdoJBLc3Ng39xCQD
J5KBfN0vke64cyk6ZVf5QKArkBKZnWR0VX95u6RK60Yq5QtPNx9fvJrwjaNXL4gyQ45b7S5zi8pk
7jEk134tRI+a9shpP+FA4mB7B0BmNPF2zCDB3LdhOY4Lp4W3QlHAh45B353cn0XqCdeSFh1wIDHF
uoIrMIaM18EwZ4+ob8JEZdLJjWkRLIjyM+hXJMLioudjiQ98ik45CC1nCGjplfnTDjH9L9EmELVQ
Z5ZQxXJ4NkadYeOr2JG8mIMNBC3bneLTnEZ8Xbmmpwvt6rgeC4qh2T2VBPtPBokA39Z4n6Md7oZO
CwCqMdNkVAzNmFyS/Hnu/Ea1FAG+jCiDs5Yy8dlOG/9v8phsZ51xthU99aUGY6K4ZZMLTDNt+Hnj
A0LxU8xX5+CLdjQRfDVZlvsR8QqA6rRUsKMysuKt1/mYU8nwaFNnr1sfTjafpvJDUtcQrXdJQrw+
XLgxmREp3tlBqJAb7XU56dU9Ka38Li4k6ZQCWCS3Dg/cg7fDtc8/t5bimp+T9o3jcBkLM1OIFPrS
Gwzr1RhTezssJZ0ZtWFKYZlP2gOEXq5/81e9dyQzVTuVZ7UIEqUYS631WyTvvLoqQVjy6PzbQ0I8
XC65NY+/I0t4+sUXI9HzVC4GDseAs2to9bLm39w12d0VUgAnqf/eosi+NHU07HfLmdc41DRIVu/4
vs78NnwGKs+3oa/CnO/o43xdrYQWdhST31ICyWlqXU+XL1XyP7Y/WDlyzi9zk9pq5iC905IQxgoU
6rhnsPcp1w21HK/d99Dz5nNPbKBpekSULpkAtj3vgZ19JCF1GDZeuUeTQ+vJs/0E4amHNMxV0dtD
yKvpdH9NzvX3YFjujY1iiiuslh6rQzr4WKAgtTgCQJqLNFK43LLcZiERmch7eEEUd6PZHv41azcP
DaknVHucumS7NaGUU8d15PC4bFXhVIKz5AleXvlyh0fDgChpY2w/cV0BKgLfRBUupovEXPPZ+BQl
wQNc0hmErCuCyU/jOgn4HpzmBq/0kpKZ0TUJZLSeWW6kwFD9K1z1ol6udps3KEUv9wG9g8WocEdf
ty2qdrZ9qq4zkihGr43Bxp1AbPR7Z1zPimD8cV+FdEBzK7VVmDliFziH8rhRF9XXRz0bLJFKQbsY
bU5hYhnnjAeDJyR0/OTciB1i4weIuiDOuGeZQaHFSueundJve8bmg0n35/bUqMAR4MrlD+P3oYe7
8aBAZ9YLGzda9nwOpWL7KZ/hUr9iktVhjaza7Y7Xmx90fCqQS7oEZ9gOjB4xyynLdHk8oC7/IWjP
z30u3zNcpL/uH7uRBBzQZMJN0T02FhQccRUdcqyyXYJs82BNWY+UHh6wMgVIrYERlHt6cbyyjnWP
qL8RwXcQ+tQjIhvrIOSqj3fkS4XLcpzJMAIpJiQCstO/7I7gbLBUoNAj3NUHqwySFN9s/3H6JrMA
9LFRYhHXaJLyHt8BnU28kaZo2rqnVIkFoy9an6htgBMyRIr8ufzYZOPaN7yMpFcLoTceO0Jd43E1
FFmXimKEKav2JOWwuqhDTRmBSfdMrDRDQyx646CHpeCvD3mgygO6n1ogHk0VjDjTGosLUvrzi8/j
eHRBTLgVPM0Xb/gLZJ+kQfwkXjbdN3PpdfiW21M5z6rwFJg0Rd0gaNd5v79yxWY/e+5LZcuLQAZ4
bTvJa1BhBdTEAdBKsmyQjNqCtgfQBU0O+Rbttc3k6acfIIKkl4jhoGsU7p2ocDfKFrjqsN7uTxxm
Ikyt+xx5TzMHW5eMg0hecPVKCFTXUHr2BG6Ttlbm4oNpQRyexjsLyJ+NvFYrYXk4gXzKUIZe/Ive
BfpeAAk6H0eyujfqLCmEfJHRJoWD8An1D5iCKzPAzxRVKeynBAcYMLvwADbYUhYfho+cKbA702kx
Too2hG85H4qneIVhLy5RMpGniuhyxXmHzGLhE7fjYlk+/7kjQdIMEScV85LPB6eMaQl0Z6C6Ktmf
VQvSBZo/6aYXEzFIyyZa9k7s5LEtdCd2orNgYGPeAQTDTGDW7cdTNb4Xev4WmxQtrT2Ozj68ECfg
8l7MJu6sZ7+mLtHQMuVv8C1y8+Hf/STvmpf3vcJZq3sHTmAw5RcbnQXM/MaMH/EqnZIBxYic3BNp
2VpFPrG3zHvc8krdMu/dwSuQ1eMoKWD5xNAh8cw6yASzj7ZJ2JhSk9JvIBqVxyoEO1/5N/pIRSy3
ye71Q1WklSMAWXcD/a8mY5Dl/BJhDNmHenzoqU5f5KzoXtYbpkPoPhi2Pxes6Un2j/ho6ab/lQib
8kCXDvf7v0Ek9ocGjHgBAx+Y36oL68oFypK6Ao5WpERHZ2gZpP/sxFRMvlMb3Yz4Hci2egdmxK2S
rVlBNSG7xcdYOqAbFzd1GuL+140h1Vf94UOxeLpem2rrEqZNiV/sXI6P+eB9zntFVPBHLW1KKFWB
B6L0HZuzxmgqs/w0kGRd8rVfgGfKxbAyOUpmz7MR9Jc19HfT9GMI9C3K8814lX66iJjsdPny6Z+e
EOUk8+TR8GIQGWYxw73xlueaO5glhaEpwFg9z2O7bnsYpMzgdQNs+LrtRjtweH9An7M6C+fKRucz
kNjwMf2CuGCL8dPQzLxKgBRy5LBKIaBUKlyleO+GLl8LWBN7ck7JElIGQzgGQ8LxKNkjWNgdfq6u
9tPCCpZsE26+WhTggVGjrza20YI7wDTPgDxNS08b3BVGcJufDivm/V1qqA0TrDPkzAfJFSeCEgPX
NnYkiUaipzJRiqASi5WWMb7HhqIfGvt83V4qIT06KF730q2TqPXXMH4urWavd4Jyezt/xMrIWNTe
9j2Z5mSHnDKXaGtGnB/2b4wQsZ2Zo7xpbl3jzT+/jB8pPsiWhOSBLNHZHelwZ9bHnizQ3MvvJsCA
M60cFn53X3tAHQPDVXzGXgrl+77z0K9Y/dzAv8CYCC27kFAHyy2mSKqFNKTSd+ZRWcCqPNfBIV3v
AU13oMFDSZlfsG+dO89GhbMSIMhMCCL+taKSbkZbiL6LqFRC+lSwUnAZaXjjOIhboGEMpJ95pGnQ
BhWId2Bu0LfaWM+c2Zekyiabb2kS3gzpSS9n1gjafJY0KeaB1W+N3t0t7kz7QOqJTTpkE/NTUFjT
LFAN2ZMj/ZDV53XQ2yMx+HaOlRUW6p0fxdD00H7eCrX8IDhVd8Y/cBZ506vjERDjONUYkC3t3w9K
GtWZiaBXN8aWlw6eyPqe+XrKABlNBp2dgyQ5nXS0TDaX+AyGU/hF+rBca980iWTrMn+c39Uuv7Xb
eTEyaHZqLT3AQYlESd+TmOl7wSPn6VKf1Wd+qCHTQ1c1KncO0APvTBG6mrQpN7gZNLiqxc62/2VX
TaldHYvEAVJX+uFqWN1F6RU2PWkqEXmLCBNIa3X2+ajtNM9TmtBQmk5OtA+S6C4mpiT3dU1zt/PD
8XIXRkS67xeR5X11aZEFfcYZ8rHX+/IBdS1nz3FikhfzMbeE6Ck6+rT8qXpJeRK4dBrA+jfsPlRV
2lPi0az9YpaEw5xxnUK+G8RPZhcjGYOM/qFBypSh7K7TyO98EZXWXlROIhl1DX5zti4DsmBYs5pt
lgwXFupFd/P7cClk8QMCEfP74LmNF1+kuU2RqYv4Y179coEXV8QPfBlM4Hm6g6DihqL4O25AnjdC
hYynhdS5Yd6O432Mw3/BNUEmK1KUiyV//xN0t74QAI/T92l/fVkUgqWCZ+uw5lQ/WSUUmmIytbsH
HRp7R+rT6Bz2VW+tArxm+7tCAOi4DcbbEQiTOWXg9jD2wstZpPAxXx9kj6OfKqytI1NIursPb0d5
Fd6bd3BEQruj6/Soe0w5npJwIDtXRrvged2DiAMpPLRlja9Bnb8dleXU22aS3JI5XUdeW3uDavDr
glI6mqOyUJ3aZOVYDosND4TJ9fWMW/sbjGwmI/5OV4vDGAK/P9BdsNvE22Ip5m3thp0rOE66vhTL
2YRaJnh3IfZ3ZL7B1ReP8u9ti2ONakI/C+0jki7BTLh/yvFj3tsi5bmPTGARVTYEvB5ghi3MfthE
2rEIY3Fnsq85+wZ/rKm8hRoIl+bDko/8/o8DkdBZaK51sdrG896Z9hMFiYeqPUdeHdTseTh1aT9Z
ihFy7/GmUsfRSMBc0kfKMwQhgQxPMB9ETq0wGHF442WOi6AUmIzDyf8ZlYjQ95kGn27aXMFXi5NY
Hx26PfqfkDeXitxgcTiqgNSVt1fNpnUHLbx1MS2a5J8rekR5KGI1Cirh+PzhF5FAl9429huXG2CP
+CrVb8ooFTnc6oB+J+ggmiNpX4GiENj6jHZJX/FW+IZ/TxBo6oDuhG0mrHzszCDnLq1f61BYiUJj
kKhZTmpyyl1oQVzXWATvO/ipq2DFuDEuzZFCRjUG2EnEvOsTXOMNNMVrkw7afZ/wNfMeX5T4k+4E
Qb16atnDhEEreJwaU9SfA8zWWUC+LB1QFt9upm5p14VG9hXM9H64Sw6VB1TyGX/7plH3NZtFButi
dce9dAw+yMRoqi+Ka8LmxOr2Cn6bE7YgMc1vTf+DeQOGBhOvZoWngUKbRQVqCucnDxLN0aIl2iqf
jN6m/4//+RxgwLcaIZvpOruSBtLwiv+GPNNOWOUmOVHXHROWz2nHj7tzDV+3wn8StDwDs8fXF/IR
8XL8UV7PK++hghrcXMyxJE8oytL7Ajc1Tf2ut+NXMCjVXzEZCuVWW5V8ZIri5z10T6txbHpVjbcq
BpcX2GDjJ6H/A41/WGwFYIegr4Qo49Su6cpmp8SgFjr3/DwVyUoj/Ok4BivfTy7/igNhA+k4nM6C
CcJzztFVNlpBGa5H8i9T2RqhrtCcrSK8bVBFdmVjWFL0QpvDMggkItHhl0JgVp3q+YSpmQ7nBJ57
owrDQnzTILWWuPAeT0MBLjtNqYWhxwkZwR7zgtZYAjX0XD1z+MbRXbvdJ1wa2E9qjNUUUYpsPexV
gqW7FIcWFOEAk3jnP6DBXzg+o6hpj84z4OMdxC5xnUPcMQjyBNab9nHP6hMFeG8GTW+SYIKz8mH+
5z672llcCMg19N0Du3MSaqW09OLf1DXBbVOcWqLqleBVJPpWLA3QU/H984FTbwEmKyss1nG1XRPk
WgAbbgchJk996iI4edDrsW4pblK6wcFEiNDbkg4/7JAEmL+xX4sUDbvtgJSagelevVYqWfIU4BPR
OsR5qRkc99eTq/pdTgQhM3Upg5jdoZar7tfBqo73PLldBYpX4ee6zfNe4WyC2++98iAauJTQNzac
+5K0ji+YUxvFT210AwpnYKC7JAN7UrJgrJiX/3Q8Pf/vWd5oLse20hySnnnxd5ZWk/w85anAtrNS
xcLLYmMCh+FVav06z7P7Ss+QuM1iHe4ywzl0E5Qprw6IOWHmqMNNHrxgfBqaKZa+l3fD17J3AkhF
fxnnrJcQw+SUVAHtLmhFDPMfwcP8fnA0GUO/RUwTvsZNCVnz3bsnll6S0pWIPjf3s5rgQ6iyWuGm
W3r6hGiDNOliu6yulN0Umd2nqVolyP6tsVyKcyISJNQBhbZmzNlkjtO0L1Vbpgl2rCSdsC7Vp7uE
LV/2lYDwgsWE3nRw++kHVLEJC0u6EH/V46nqRuRxNLRjjc9nWFNKWMvXQ8FMB90yjR+gte466WqX
/OfLWK154KnOHkDxHv+1XvnQ20gMgj7rTocV0Vv3yXhaVz79kN/TLPOJYw0Fd2S6f+ixm9dO79l9
XnmKdbqgmT0ymjTkgZK9b/75m+P2qf4hL7BHSk/rgUW2LaTSTXbkw4mlOCBMwdVRJyEcANGoMdat
9YStpgLSCEWFayIw6Wb3h5Jmyu70SHnGsxaDSZhSKMvV/v9HVeKIyCYdC3Q7u6D77tHuI+smWVXT
F2kWz0V/MRXjWPLSdAp8SJLnP/PUc2iCJegRkSx8qIEUuP/T0dIp/R6zsXeAY6s6+Mm3CcyKGD8a
qLDfGQWgsZ8sERlrb4q5c87ZxUqKkvmhz28WxxUWi9l97hwXlrdFCUpnXUcKRVZgz4SuGKWe+dXY
HNtRyMDoKsRjbWAw2RPHLe7XLq4mVwQ8oSZz61KHuO7oOt66j8osMBkNLfkmJpHl+aNyRMa7mPrO
ypDES88/dpXgfsqQ7BHF6CZXXTDWz8wkhta1UdPoyCoL35vhrVyC6WAwQHiWRXL8JvSrpke6rzXb
1gcRSvMQ1DD3P/StEqRQ13KNUXJJbm2EHAYGMUD4OXwgyHFmaZ6OF7SBzbfRlFX+JVNNG8u6HL+3
HFMf0xEuJZAXVyhjTNNI4znweNZrU3wc9WKc8U29pxROZrEpajzXxgCdAIChBdkUM/+AznIM3mkO
9nnhp/nPSs6A+eYsMhKaOF1gF7u1Jx0GraLysycn27XYCaiTnhumNdpTHp8X8LcJNqXmdcSvVO1N
xmE6avLkNmb+ZcqIIkW12/trNNKNpnOO0qzkS9OBdDgrJy4RQ1KYYtUEsEqtvZKbwhM1rDEc+QwO
pOwJmPawzX+0mrQnF0H1vomVJ+uvkb6mJ6fQW94lEgZy/isMSYBSIML5d8pRyWYl+bcA02KEnasA
leIzHtmZ1D0mg+S4r0//8IEp12OC0xbgIgft+VZqqnlNQDZDyPNnd7BzKtNw88n+l+opqG+AOSj5
iDJHwWoTIOkwrgo94Jpieb1j1AqKySdxvpRT2RvGvBslsnoLTCx1Gz3izXd4xVQoHdxzXdrRIHfD
NnpRPYNCgrz5CI5JuMIFYeDf503hTQHOEF8QgaKwHCBaa6AXs/kBcGcvHFV1T5DCKPEmFLUC4I74
Lxl9XGjErON3LpC/Z94xmbd73052/LQoXsXTQG3oRdXj6eGDBSzrXcGFKhVnwERBYlI29E0WKeAV
AZM5ReWYidsO6Rz0IlTnq4nDEEs/qrnZRoLofKHUxxYEK4RPIaTQsowm47llYN//jmK488ChzF7C
OPmgaTfNwuEBlRK9xibioFV8dPfulZj8vqBVoSld1UvUd4D8NUFK4ajlil00TXWxgDJHVyhaTYpZ
pqWbk9xhJCfy6/tDa/ox58F5CRljGS+21it5Wrtz8a74fKe0BDlOkPk6L+ieUFGi7iBgiP+5odo+
Ptw+PruuwOOoJ8RHaGG8OWJZetcugEDv0FD9NZ10y7GENXkkOLAAHD+J2mLHG/iz6pBbmGkLg2CX
aCDXWAUQcL5mL8MYZicpe/3ExgZsaf7/bz+Ps4oQ0nR3SJQBE3aiZ5qI9J4yCNp9xpgjBB8Tsw63
m37r71YQlPzuWAWEuWJinKDIiyK91tni7V7Mvk7BiBWVYqMhr6P09tyvOxRWy7dttkA4eUC8l7Xy
HLyJJhOklKp6vtzabyLusGHV5htNvUWPWfSSnxN6XNHlLRlHwZIn8Zved9CK0JPv0OZfhgmVJXJk
2I+EVQ/eWFL0zG6r3U1czKM46PrNdLRK2TBFNVp8L8pfzkw7FD7eXPuQpO1c3FNeM/5XDb+DE2jM
mJkdBxN6uD7IaTtgVqhjK4BW82bMVflgo/Mb8966gdKhws9cZuXSKxKrIUs9Ya1yk1Z2RGNhLscH
AvcoJDjomRwF1uj9q1tPfw+gKRtSqmyu8B7d+8O7vq351oD2B+nOzgMBQZ4Xmupg5G/JmkQ/l6av
YEa5c/nZ8c8JBVOdxKienGBBRgSdPErgJ0eE1GuPBppFaNxI85wvGc+6Fyqi6ZHgQVg8gBryzqti
ViUZv+W2e6y00sRcwnZSZI/gt/Bi9wXJ+m/xNXvrnObFaa3i01scE8+uVgcn8RnUoghfqg5hqjEi
fybIzR3vnGniy+RQGpiXkKYGT29UFXhooTtENtpuzukQ1ZeEUAkSEO4pXp7DWJV+PTpAmlcgQmW+
eZfYXm6MNzkQI3hgSpe7Cfl6E6QwohIKAiVWa8L3Nxv1kFos5o0g4r9PTlZQvA77I6p54SNjC/0C
HT9Wy8grsnRx2JLLjAYFiqbvDZORR9OkAAM7L6SDokUNXDzlE4DoV+jmB0hnJlxS0huV9IjBwmcW
AujED2DYOsD3IUXqV9uEaW444ayLVIQc+YoVLXtHsgjFR1RNwyx504/o2DX1qV/73kvqPwsUpDp6
IG5sBpxN2rS+RoCA0LtP9SI2v3S25QztvVr+PmtM7zO+vc2IVT9jZeXD42upKdVZ8ci8irNrnqNV
p7d98e/16G3lClXLuSxheTMjp4IUh2+v2FlgbD6K7Egd/xwLnY5s+xxjnpEoO91IRMKiSpiUNDJf
cbDtUyDqEPJsqEZxxWZQ04acoSBLGP7cBDsvL7PM5aPo2R5K178621QbcXpAB4mu/xxh+gXdgdH7
tJvvChXxZa3sxSE9Zvxe+kvz8yY4m+Z1jMPzDMUrSueHrWaQ6JWC+JazaVAlRWlhe1LYLlqnMrGE
kGYUMY9LvOb+X05A3LKZ/UDPwM2Rx8WADrGe/uWEs8iHGYFgfJnOVFfj4KMNi7hHHPJSlgw+Ruls
9Lf1lGKQ5A9BgEiyfm6Q/dxC9rE+DwjcKsHHOHZCDgxcmDiqO2x1VQ3UJSisFNAhmdRNFrVVjYmT
6V/UrNZkYE8OcPaj996thXnkS5tMcu7s3GdWn9oCSRtV4uvVKJLoJqAgX/DfsY6I4uPvOdJufoDS
oUO6t9ReVdfUa3zWZ2OhFURYzKTkLE6VBHSbRq4tHf7SgOHENtEyooUJdcszZUny09Y6RBQNZF/w
VuRyfar1UDLxQZVyNxYlcO8tOafPapmppNAE/k0WqeoaS0UgQgG6tYdsfcPuStPgFBE+EjtILHqy
fpX5HEJ4teUG+euOWj4nm9nye82258oh7rtlFbTbn4ja+/EoIa8VwpmlEj5IJe1jjzL1XdzWQtIo
iR8NhN5lXMhg0LAZVVbX0+D2ZjVuHqz+89nVwosJ9O3wEbsJJRFPQAlXgf7BUL6kx0yJnEYy8iew
RKt+VAn8+vM+nmuxW9SOg5SgCV9qCp84pEU70mnV4CjA9EU5wSFDAiFafEDuV2eCbo7pdC3bywjv
+4anQCRPjwpfPXJCTcR1O0Ic/RNqB+OsXnTojKvzu4/BgCubxUDm4ZvoXFyqS1WcLP/0707hJfFb
V5J50whgDTcCEsnfTbeCRrtQ7WzWEYhRmKqQaLrKhwvdRBr4+TXK1q7t8U6p7hb5notee6K6SO5L
iSKlNcyFomIv0yVhSgG/LkR9c2PVp5HXpbZJVSgU97nu6n7Piwn4H648dRb8ZrPN7s3miv3t3mPR
ACxl7ASMqlyDQxxkuU2KlBv5m4SVNb+urPQhNBM2JLM+nr2wf6czb3MWc6Z91ila3mUDJsPtqG9o
5vvrAd4maLF/0XgiziaVgKRyPzKfN+MzRRI9S+jLbxtMVGMYTXV8eyy3O3zeHntD7JZLD42VVD2p
v79DHCpbFfH37cSmmL24YUYieZLe2ehhwrP/4Wmm0Rl0YH1gv0JCXrhWNPnTAEubfxFgiyggE7x0
1sqEntP7XIpW8AjM5gzzEkZm7jvDJsbujngPxBkzyXyMyXCaD/peOdw2eEk9065e+Sca9WpK4Ufc
5Yv75WriJ36W/qD19+k1ZyRHpjr/6LqYOsRWNw9DylydG9v4ImNCAyjlmBYAEHaZfs6m+h+8GROK
lXXU81obkI/yQx/eimS9jGyc7pAJIpmLAdCew+uxdEuTiiXyKdaCjHONrTdu4mdVARyeKur/200w
dgOZqvUiJHlsEOkqwLcSI4fjnFmypg47wN8Qktb9fdqKRunO9BXXpe4iTmMnt9esuUuzlxXoB36y
q/nEkh4hYzueAnhb+4FXZz7FRwFX8uwBwuqquVdGVLYA3sQhzl4HPHluZRNAHv7f+SEjvM1byDrR
8+gOBhLreYtXb2LbGV5YtaxF8Io6Y5+scvgchhJIajFnVXIhbys4K8OuXJNkQvuVefgJ77dI2U0L
EFbsWyG6bx4qJLp63NnN3LgdTTcyGE4gagtjRv54z931i/OF9YHr23Y9XzDBONcym3WddmYLragS
/FGSUyNMGgdLSMuz56aEvsf1cXbXwDtYuVxSGpYC5FSb9CFZkGhaik6SbFH1QzyKw2UyrkQTAUNs
j2+2OAMVH6YEWrFytO9rgjCWsPNOFsHaEqidCHVXJYJQI/EmxAUJpqChP5PRxZOtmdB2aMkMdwrH
OM89Lk3iw62DzgSyrWaEyN1xc4RLdp2+JPqExIia/id2t5NJJ+hazj5gLYQqyMKC2hi93mL8Lyv1
o/IVXDWBhxL70+3WRZYUfGmeF5sgq3csq8RcoDAOtYBhVdQXTogsxRJjuCosO2IAG4IFC06nFruL
kP7hIb5AQSZWsGE4YGcHzIhXFYYxNAtWHctmoFv1ZH4RJwJBKJNnlrUbv8EfTEFndh8k96McMl9l
B8+loBgf19k2F4F7w8bUJHaAKlyqFgBDKV0W5X3G/IT2Gl4J9OKnxuxM1rvwJjeiHkXW8B9+fSPV
PGr4+sZslEQfQ5xX8uPH+MgbQJv2u5dzpUsAsKOhF4pNhKmZw+pDVJ7C3cY4fN4uBWQBil9bL9lo
OgX2MaTEOyhsIywoQr/2LiGhjsL+mpujw594yptKXNIx9ZA6zMd0o3pT55UWzotvLRibaAa/mfHG
mXJlfxctYiX06C+yr35t9Kq+zzx+9DljayxELSIrwD425QLutFX0BuDs2Yv2ypjqpUCP6E0pdnFH
5nVNQ4dOVx8PXo5QBu/42wNDaBD24t08RszpqwncZRr3nX+Tzn+pLzaBxsmnY7r9CIEaTiEmp016
4CTEAcxsFe6psMiKrFrCbBXYxhCGDTbpEDszVPJ2rAUbBDyK1Lh/Qkh4Vr1scNIH741QZfeyumJx
lnm2VHJ76QSjJZR07DO0GJLpD90P0AJFDGaLcndGPy+1sOs+aR8O4o5jJZlUTVGfq8Woi+AxpD5H
bBA3mzkBZfoTtR2YV4J1GVr8TIzm3fRirh1G8ihozf7kgKyzRZ8S3z6fhR8n3/mmZ+/V7x4rrYUg
SYWsUWJdk4oNDJ+IoB2KJjRPtNsv6TGDNaKfSovz+gPhpNpQW2PyYnf+oOR69A2vxO/vBM5RjTxm
dhCzoyE1NU2bW5rWZ20E/xLLsn2SP2O/L+3DAaIq2dByTxw4rnhzkKZbkSblRSLNlM7+laGPm0N6
rRreUMdrcAQOeJsV5fnksF/q4ioep/zRbPlFuOIZy0mRF4BM+s9PtHaDmpM/yvMchV4NgZE4CCDt
IbOGlgiuTmV+Ty6u7tOjRPUC+13tW4iLYLMwMZv8Fw3Lu4KxA0+QN3w2iVHK+03K5UktmR/BO92M
yXbJEnjjjCQsO2tq5FGwqbg9sclPB8lkm1p8hqDQDfUeKNTQi/wwuNDF3XmKv90nx1DnRsWxVfEf
0H8QjH0qaMKcT5NhOcJNFqXFZ0eqpMOj4uwnlhXiwrTY3ug49m9Z78mimmWdPzlSl1HUm9HAF9oL
12IJqRr+6QgJmkYtxfs9onotKnD15/07t4p35keTJVwL0na/3AhsAPkHsnwLBtHNyqSvAqvHrUSZ
SDhWlhLxsOYBwLmV8EJt8kzKEGmGY2SMzlE5alSAcu3fLrN6RStMhF/AKh4kKUDtXygiHGkmErOG
9W8APLtUiA0b02zXmsygKHlvjXH9GUbw04BT5IYAncFYfeotP2+STp6xgpfRMA00BzZ5XYhMHZkT
6v7k3/KRt3gZfaLqI4+s8LKMIC/4Vgiv858Ag+ANYB9d/OMTwnXUdz5GEpeU/KfRDMR7NzE40z5h
KWtYuc5pQkRJVpS9zl+YVkI5LcAmy9IdGGz7iZ9LhQIx/qbd4eOq1neEirDLNCMSRYyBbVTXCoD7
XZsggkivC+8zHe4A7Bu/1GMKkkyZcmfqpJHyyt1aQYNJR3JQLyVUbUb4ssG+EPfug2d/uyOdWLsO
dufAChgxHQZmnVOpJnNtSXfz2pthHgQFUvkvQ5yAex0C9F3dYWBwT+GykWMHRl6wb7uGXbSHV8Gn
Uwz35jp6n39KU7YHvl2tKOg1ZXWhmicrYfJxgRrcg+QnyIAKN8Pz/ONk7WRH1HdUtROW80GVh4Mp
2KAVXVDLCRNpy8FRz5yJNOct+0I2n4SGWrwTMF1A5MaqjYqqzOZIOaKoFGkifFVKTzXTQAXNpTUQ
MiCNaIytwrEzV+8psxxk/PDZH8Wi2jtiOb3z5CRH7Vu4fi45h6ksqb4ZjmPnB0FshtL7mG5fun1M
LPfe1baRAtnB7aXqWmAkA7L3jmVv19bqYTNpwOn5XoYRPP4yqP2qN8ULkeokPrNF1aezv1GT8RjF
n8WK+ujJSUPtt/Lvd7d9GtJBSLaXMdI+fA515YT9PxrXaxgmWMQkyk7YDZ22IylO/FMejyLRdxRJ
A6lRkgWPDlbN6P//Ab+W0SdQgguNtemPAziE5qZtl0PiTtdKsCNAn8m0NAlBxZXP3IhFTSMoRuS0
pmhHb7rA4P0zxaioph5nZPLmPMqgJ/aAa8mc2Biut207RrX1yOB+rQhIljpSrrpdlqCJkfSFGo31
VlTdYbUIJJMNRJFvi0TCyClJoGIlInfpPkeUBhkMGT5pgrz7V2evsNis2wrJI+y2b7Le92JZUNXW
HIU/jUu2LY2LPIE41Mp5ByCaEhLM3p9AOO9usEsWveRYQvu8ZdWGtMIrIZAb43ilVYvPPX6Ie7ab
UEKrvAZJ3DDAsqoArJX+zoSDBQEKWpqe12uGk2dNM9eeRQH/2Qf9mVsSYh0AO9CNDPlge6aNaQ+K
zIYpgBqYpvBdSXEUNZS9u9KQV7YzszQF9S0GJeF7ng5vD6N09zVjtPtu1rxBey28LAAYWkUMOMLG
iFlvyQRExrv6sqAWD1nbaULSJVphRdzRlA1Vfnes4LmUMhEDg5fIUmdjwBd/2B0vMA0GWpvs572P
HDWs87AZTpkC/Ebn5xaowCkC7jnyUqRhCO3sqolULb+JKjwP2ib/vU2G64fwupBGw8KXM6mTaI4/
Xdr8eSdP2J/Cvo3yuBy4T033398SAiG86bVmx+j8uxAvwfLoSFGpSlr+F9ttf+ZIbJetFbPdyDPq
8hHHVvzUvPFwcvA190H/cUX6wZ4LzZXxyLSnvCoD29aA/dE1+Gf9bA2xgO1HeAPU+cGMUK9NF4v7
qhTMwPQl9LzmgvfMztE5g8HPe5ytT8V08uqB16geBeq/xTb/1OVQxXCTZGEqVeCBYoNvrnH1aNeM
2i4FKWTI/kfMoYiVd+1qJED6+MFaAOKVgYid9n9kW1twrVlhGv/xr+3iHxfEnoaMhE6M/NxLS8OF
GA2Rj+uNnAj69WefscRniZRZW3rhu8UmRIHbCyfikG2IZM9ETp8BNNYS3uKXTNniNpeqobusMnjU
3GGnYFL5JU+tO8WMhF1xk36a2KBfwhMCkTabTIoL1AVdvFo2HooDmZHSz9jWAaj7tUFucqRzOk6r
imAhfvOABinLHdea36hOursxKc2i/FGVM9fEBEKQwrqKX4+5hv/LsfxuUknj5lGR5ycr43HYcNEk
4TJ5ey357Sr8AiRDbZnsXP20em13SsV7rUZsCNiQRKwLlIn1ZbzSCbYxiql0yDzxxNVAGsCiHA/a
TizuCNm49BlWmi+1+V/G6VtxhscwzQZCvmmo+/oBV4v9ZDlDqh0mn6r10c6meWmvrmafQ/wDpnHA
VK3522e+D3H9tc94lySx7R4AkW/iuYALvE80P1diWcZW7zKziMdMhWMckN+nyBLKcXA/g6AB0sdi
QuzsvEU9cHK5LtPZQTV3wehtXbm97UEFDjMVBN1Vg2q6VLBQJDcKRDr+0UIJeBgEyIqakfCfly31
owlI2DXwiP7rSspsSRE5cxEOIwAEV4b8p8ByFCi1dQ1hSP0vBZVO6cUhuSnHycAU8BS1R9vuizHG
W+9VLnBEEpRMi5cxKlz3DaJoTD/JblTBSZwdMnY0aQKgPCXQ06gf6rhG2q5ROf4K1sAjcyBvgJMd
dINAu6LJJE3zRAlmXT4Cx9ltTX5n50JpTl4/G1jcm0i8fqAwj5ydt0RpiqIB5NwA0YTCXnB8Iw5/
WKDCPxotfvobx2MFlZof3nnjowERjKfG4lOp3HLjWLVErsranJNE6qPWOJi1dE+LYp1HKKyvAgsh
2fgGlp0mT3JF9CxW+VzgcjVZyeBUTlUdIjf2b5VLnTaZ0mLJTN8NX08G+uSXr57QBRUpC06jjZt6
c5WW8X0E8/ZwrBVz6ab3OYRXgD6omX3jXwEOf06Gp/R4hiaZ0C1weGUrWqHHbhDbjhD3+nRmK4y/
lpQ47ibxowmA/jnQNzDyb4ek5kDkeU+U1gYSeUSYZLR3NZTZBeUH1rzFJZKBCjpM8mpOJYctsZzP
IABXtWmES5WuwvSFJ451k+SRevrPw4UchMiGVEf/+lm7Ij75sa9vnJHw/mKQFNzppXaycdK4L8tr
LleSPoS3GgnwsQgEwPVYBjBI31FK9s0mKg1uXBrlU42Y9CRhL0O8dSX7mA24P9U38ZnadrtohOZa
cMxGYcvRqlrRH3RBh8a0/vzk6mALTuvoYDn0JdTKko6YxynR06TQACTQIojKLfxC9o5Sbi5tM1WL
IR6wpcEe9ezOphVek75o0td+YyTs+SI5mNNSifIbr+y1LDHhxorC+EkbdNA5YzQ/B51979cEVWHC
a28bgsJPHx6RzkNj4EC2GaPcyFxr6qMjArj+jrelzPMf9ELJn5Cc8RqJADgElLFE8/qld4k4S3QB
deqVb/5WUM8KvIGRiTMyXm0ryQk4I6CATsXXW0GinbEHfeuAutO/6p9oG1VCkHQnsAZ7q1LuPZSn
SoEb0cqV8lNuBOevuKC5QIhWHzTOlt+aXAnzl11MBNqGuicBT+p0QJC+q4uxSG3mex3kazqm/e4Z
0LB+qHrwwcPAfRpBVyIVQZCBRjljeHPK0dYlPcI5Ad1BuaEJuZswtzuR3KaF01ysCxYGlvZ96qEO
4HPolxe9cbeu7xNEj2sW1LKeJSg3ICcUgJcF2TQUwZYPHDBfFlusBQeh/VEvy4z02mME8cHIrC+l
PR9GEg2GAsyN1kYZC4GOKDjYlzTQZnV4hX2ONLHpjk7krEh5Y5MB5e9BTGgebN6O0/UQJRYi4Eoa
P+oaqRXYBizKeSU2K8Ugse+mc1qKP3BnyAuyXvinasDtWW902zymUAeIeG4jwjTGx5k0rFjNkggr
CbdY+xlbbb+vWP//tZ9NRj+C7BzEt84MQMYcNfHyWIH7uxQFbFujCA6Wm5kBYfWVKHSl7jwwBq0V
XwgKUg997pk7koumnKl0TVkBstX58ohddGTvZfgSE/2umm+Qk4sVxjMrZEGzhsO9M2v+F7Ot/XJw
2oweAH21YkpePoTbKwGEnTcEhhw6tGazukuRtnMcQpAdrvXv4ck+3+XBdRC/LnxSaRnz6Llij0/u
Qy6u2Y8kaAZiCeED4jUsUjUvWaPh/6tYHeU5g/YgF5NKjK5hoktzX42TEIUNdimgtbz7LeD/dgjR
XZNIAvTwoulLfFGrOqOlV5q2OpLKIaO8/Pg8ZTxTyNpl4OHnpXYrtVoH6ZWi1lYjLcGx0FAOqW18
e1tX9aXOK9MssLlqtSGoQo2kDVkK/8Av8M/LD7J695zuXTBs+TnNWAKfqSZUU79FUMCuRRmkxbai
drvunnTiQpCQ5i7vyUaUfCHYlGCxKjbrzzHjGKJ4uJQqKK9PIpnmfO3YjeD0C8NcbK0mWRxFoHfD
Ebmc9d/wjHXrDd/T1rJ2zXJvqYyEMiKydouvCSGyx4l/nbbEWFJwWtaFlaIH3T6LXpr+HEMyGW5L
jlPv87EFHvcigdG2wbElHETaP8qge9FQ+kU3D+Q9gykIMifiMo2KiiJPiqgDQZIKwYlY+v2g1dNZ
ohG5kXx1VH1ADOEJGS2p0UtsvYjl8cbqFfU6wpeERZOdN0JbWlu8SF3SqVE8wQbJG9jLQO5yVV8n
2k8mBbySdqHry7V0SSNQQpdwD3T5nL3LV6IxZTC6gdDgNiKAoCTckjRNLdtnCB46bhfvUbLVoHf8
bxalsF/MY1gNCNIiW9l4Z4XZdS5RaD5ZmkUfO27q5Exl95nw5qlYqHXk07VC+oalT8QLcLf/1D+S
jfKopl22Pr1k1+W72fUyDyVZJmFI2kHtj25dRDw3o9jCGOVor2KTjq5Rj5VN7DH5IFDvISD3BmRn
SQWw4O6D17c8zjTXt5jpUPi+L3NZyHltNh6GY/5n6pfxPpH2WzOA/AxyM2M4O7V6f0V1WQoQsLQN
fV8JxIL9U1NvRIDGqnV7vBNLiL/7bTEZM2lStiPgJiXd3E7CYRm4sLbKBT8pFRR9407Zrec3Juwy
Wo1KmaxZJxHPIDwT4DjfN+QrJpUvCxA3+PZxx9saGBHkPX6/hVgkzwuE/XqpsIeHRyew32v7Uqo6
QafI3R4p3d8BnhMUWJJNZmYYrwXiUU67Nrgqv24JDOAC6y+jHZrUM+X0TO/VB+hNS8/jpqHbUYhE
GXmDXV1FZ+UF0mU6CxTpBhWlgxFtwCMiEWvNPUA91folvy8RnSxmcoU91FXmfVCU9UH21+yEr/7B
eGLhFXZ1g1RZcLGU8NzVcQBuncKJKOWzfx0i7Gse4nWps2UsOJJdBIlkXw2kK0IVpha6XVSLP/qZ
4BrMrtzq2/jYnSODv7mpICq71NCAFXw32c/jnt2FQ9n83RWrA/kUNlZF28Dup4xhKP0YmGMk/1nb
3G3K5I5uFsJkXEtGsEleKe71NjeTvkcJ3HxxFe75sWQVOCCjyAaEMpr9tuXO2WzM8tcb6AkIykWj
Uq5nhYuOpbcuvfF9BWdjZgXclooAr3OmFwi/aFFoj2QHAyZmOCGlXblspxXCs7aMqecjdAr3mows
uEDO+29hYcyTSulWrHEi8Vx3XDUL/KxXSyMCyJLzRAvtw/S6SBdXbRcNaDwZ/TtULc/bfnlGsPKS
rZK8nuQCOUhle25Wcmif9XZpYcWtorlikP6YulLh8rmxWCecbCNJU9OkxtdX92sYNwHCvnuDyClz
PEod8hfKyyNqF8Ec2zoJiKeMStTTinfI7cGNIoYB8pLnIqXB87KnGoKc6pUtBRbYPgOFQUk2k0R6
vC3DlqfnE5jRJLcEerxSGd+GhkqYwhIpjjD887b30TopXUy8DK2S3y6JVUMwnOWDssT9JqeLHJui
8Z8vVDYiEKqtCIIXqXCBiAxzhPp5nBUwA0EX4FmE1F6CMzb2MXT0TYsr9jt1GipA0BTLXow75nst
mUcZQZI50b/FjMb3pep7x0IqaE/6eaZfCb5L/wDEvM+rRWUj1YROh9e0Pcj7rco0K2bS+VhzIiml
Eqoj60paJ4l6LnVUc9AA3Stbtw91lYXhDk9oeahJrmHO3EP/vror9SeKoQthsHz1mvJXSalF+FCi
JkeZJHup7jyKG8lP5C6PMYwMStUnOPKGUtglwSoPaJ0ctlitWYou8Y2gQXi0FZfiVvlHzD8YPXV3
qczrepF5Q6fCCnb6z0uAwZ3qPt73jVWG1I+0IZymAWXZZ78cdXiSsPK25a5yB5Lj3x18KBQzSslP
+3lpWa/Pn/WncLGZDbqcrDTCwTFicilfRqlOdTREtc2d4kgPn502wPw/xh5+LFmnfqYwKLxLScTE
Ju/UXAosp3ApGGzb0f5CxunnqHrz5oc0FqOcKSfkTr0WzBE3KhoZ7LSoPTiN6H5jzm7RjThek3/5
+N6ynXGKsw0c5aAnJcGzt/zkqSfaGLqlhOtB7txcLdRb9l8PqJ5N4N9t3MFWR/FQ8LVeas2h3YD7
3pqyoqcRsNXc9cI61uOhR8/l+IwCKbI2Oyhs+WDMgovLzOcLBDraM3tUZwQwXP5lKS1GAjvdUXHJ
9XOYPwCy7RZC9nc0Cj9j27t3FHAt+LkILE9adTUeFZVeje5SpxgqsYtf9fHAWfKjvDva61Vll0CZ
HloL5b7mQEH7AuSjiAFN0JqYwLPnq1X7Lp1CAjVW2nAivtRVCoWzeAYYhrxRW1jmyrjocpVI8Ys0
Nwo4OBHYjFls+v1N7P1YgqybDD/hWoLRyHKr6Zbdc9jbOX1A/haaSXArD5sCRmFa0Qd1nI7bTh1s
vmNW6JwselleMl74A7eEU15XY+tofgpdMpYPydnl7sCmhgi+IhE7NXDbguAWhTizOLEc2DFkPugp
AI9c57gHLOM6tYYj49LYUXNzDNnGZdk0+iBkj7V5abNGi1CSrBbkO2BCl689rgw74pNUissajnXE
SBbicetdMrdelLM6ggLAa4Fk7zvBCCsni+fdyqFsanupUh3IFkkoJRzIfLxTX53RfS6oXtVn7h7I
m39jjHHuTWeFBSrcbOAo6VkclccwUyw/cDpdNY7xNdYwWVCL/zAgYsJdVc70uUQH01z0aPBih6cV
9g9acX7w6SM1uc1SCkodmU+DGDbLRkl1sQrS864pYFs7Fm12Md5IWpN8Vi9XYP+nwuuaf3lOUkCC
ANqsIXozWNJ0eL5g9Uf3C3lhu2UKrIFBzzkHjCpT6wDYEWfWddmuYhvt43wzY/BpHTv4mWUqoyMp
YwBZC0XqFHjKohtdp+1zZpPX70YyxtmaXRP44D3vTvmMCU3aMw6eEg9hm9l6OLnE3LUZhc/CDRMc
xm6E5GuqLb/WylFGOEV0F2zyjrC1h4bwFU5Nlks5+p/gEJFnnhU4OhJdKgXF7Ulw0+b+BP+5O44I
Wv7ldS0TExrZSrUAMl0kY2z9pTwW/p4bSKT+M/7fWDrF77ssWVKm3Rft78L0PE60Ot9fKBef7Gxz
2vpdlfrK+b5xD/2vC9GDXay9QBWdIDmnAtkJ1FqMCVQ8Wl5cNMYxf8h/da5EwWkn1oOihvkb5yBF
8Rdw2CBTSyV1Vs/67MS5xf+Y0mgqMlJ1C96SdwuQS4yK/NuhTIKrxRVsaMmBJGZCfDMep1peRlgY
f5r+0hcn0PMqiyvZYpsPw2548FMmrbhjptRlF8K2E7vVnY9erB0TGtUEDvUGpAb0lc8wuvSWi7PX
fYaH/ZgnEetLNV4q5f3yU3TQFhwafKu9R41YVFVz+x8CoSXyuWXsTMaiA5/+zDcit/pXCASlYRF1
BQ5O20p5uPpqKickR1uERl5wP+I2ngdtMRAI88mbK4wV54e22PqdT3DcPyw8qpd7h7mQUy/X7VWP
ciFHxHjKUhMRKGES8X5v/XA86CYy0sIRQ6umzPv4M3FeL0ctQIxYgQ3BYJyp2i4xg1dVXrJPz/9z
pkfI0+nQFRBEUEIi79sq1pkXjqJBBVeH2K91MkJWzQhVbxdvNB0PZ/UsXUyj3nK2Qc13g9I/S/4p
Nfuh4k/cjvM3B21jnCEY4sMi0UDd2yNvkbo72nxcCfOhWJ3OPhrSEvUdaA24wIZjlp2L9CKJpvPO
LsuaNPI3DQJoN3j3B/QQ3zF+xtgstQARn9yeJ3ytw+hry1PKDZ/UXmgazd7asLZML38xOw8Aqk0Z
xQg24UPdxjL/pWEKHnLpNQFIsww8875jeNOClJmDTtnHfL10JpnHMttk6U5lNxfYaSUyTrblQ26/
3rTtFc0121NwyZJ2fKKzr2742b1u99n7agP2bOmNsbDwmbQ72RqQFcyLod3creWIbrNJwc6f7m1m
FAz+CFRZJHOyWaczE8wJF4ue1rwTG+s1ghh3B37caB7YPMNl/gi93oj9FQgXCyNTZiFrGzXW8Omq
EEBCW151NuDpaTf4i/t8TEHsuRZ/kfNmJGYvbiLauUayYz6NY+kntRXVOJ5MKdqf58g8hA6+4154
JBKRJ5qO9ynjYLkDf7kHjXyEYwYeyUnnHb7aw17qSaW/o9aBDZV3eyh465ApyJTPEpb+Oirs140r
RRAvAniEAhCW8i+H6gqvY4CSfC0fkirLPWBMFIKwSF1nAGkMAloPUPy7mYW+IeObybn4gNl0OLVb
Vlwok53ECclhqzpWk3Hv77zLbWAWSpSnXSeyiasOK7qIpcAb/vg8AOL2N7AqB89qg+t724dDZmkY
ncXEHl9DR9H2fr3KCSFCgksP49xjEjdvx14EyWfBsbnwk6frdGmY7LNGrkHVNPnJC84sMOvox2xa
ea0if1x/zVMo6SVBWwLenTMcbz455K8c6jEM0lCEmV0srgWwolHlbAXlpmnExgPnfvvjKtM4cbHU
ZUkClssoYYYKlCYJi84SxzxwDCL4/qWVfJ7GNVQ+IliYdGyfdvMJ6rX4XImBO3x2qmKcLqiXAOJf
x5bIzipJI7nyspwAamEwu8sWRzOw3ftsVHpGsQizA4k45CRC8fswGoyNpS4sw0pGAhhoND94fUg+
UZ4KOORQmY0ztThmD0F/h7LVvPipXkflOBwnZeIWh/7Yohb/OJ1D3H3OqW+OnMoVzKg6VRJau0Z+
pCPuFL+m036ZjQawOzwKg/0I05tZfOfLg9/apmNBtBIp0ZSwv7E5rbpTFkssqnVKVO0j1Lf/8C9z
KlPaWg//AbLx791plOmu4kxYIRJ+R5iO6O6lzMloDapyaCJ2JgaLAAwfYv5N20iTbd5IEdyDLRzX
TYf8rZs6h5nSQ/RDQIcg8Oa6tw/92YnItP2RFp+yVRRtW8J2OWaLACDnXGwqkU55eAxBp8NpozvR
GEiZB3hBGP7WqsR00/OV7cQonsy75ePaRPZ0AlKNfDamifPlbq3Q8dgDgLpNoWq+mJgpxv4z9tvz
TVu1qXLCF1BVfiz9ZlR+mpYoWUMLorMmPjuaUxK/mczIyJ9By9VFGgjrh48wdhw/fWYupUFF7mOh
hi5j/qbRkd/fJY0pD7k+vvJmeD76bY8Z8hNhL7h+Nk4MqRN5miZVheJaDN1Tv7/dpiQCSi2kCjNy
LD/rAK2dzsX8hF8qV5DLaYO3IUoo4BGy2KGDMuLlt1mjoJpvX17JzZ18THAg+Q320pIk18TbivTN
nL0zCXhnPqEZhHvptoY2KxTcV+hXH3/rY4H/F9RI6EwdhN0RMKOZfZSXntBGSGeHR5YapjS6u7xC
ZWUj0qqEeBqkN0AET/COEHsAqYh6TSK0Raw/W1x8MuoSlXpuBLq0kH8KvVc57259NkzjoP2MUpa0
uzMJ7WUw5tjkKWrEMq3kswBvG8rLWCni6CzpQZcjKVFNRJeDMB9WYWW7I/J8IweQ0p7n6HCOPgUG
fXK6u6WoUVw22/HhbcCz8xohMd9Q3LaKNRzJYCjw2zSnr95fD+zCXE+7Udmw3THnxSJOXlZu4kAz
//BIS6qssryHI6jdSDasYvHjycr3xW1X2yCyoI0qs+G1av1OgAe7AAqgHqiuFRVK6/15f8f1kqKL
s163r8d0r5Iv9MblrCTlDkPWlZoPKGbZIyUrMsa6u/oXI0mnN1XPVsJbYqmlyipInrJi/lLUpHzu
6rbRSX4tF6G8G/RViB4lWpWpD7i6rcuNUV5xydJ1ry2FKjcVh1ReI2oIZ5FpF3tQ+16kQfe2YytC
swoybWPI6laRgFDrt2mFOev+xwCwO9wZCU8NsU9nn0Qezj/rERBJYUGbYZonCY9TPNplPOrIcr29
6ydFWj2RSOd7iLlSd3AmUmETar1CRU4s2VIcTyaTTfuDqjnmGo5wMoVnaoPI/jDp6m+QN4Jo0Y1O
+NJgi/YE2GS4sLvdugT+UsGsT3KlFdbMRhjLXPqoy99ZgTaMJ5/jm036LnFlNaRkvc7mNd0UKppY
f1p2NYdh1aJq9MbMdoo5MszbO7kJcm2yMPvscXE+VFrU1kAdzc3C4CLUcoIGqPAWPgtkXr6uVJI3
y+jHu11kAloudBhaGF9fXiPLOZF5t/0ZM53AHaQm9aU2ayQ+KGPdLHMDnliprivb7cwhr+nDvwh2
ELdteaAAGeN3W6QyKmZxuF89eWz7LY/Nf4jzHit7b+mgNxzCWPhodungclBhg/wxy6jd298/cOdL
y+bY1DFNmA1lFMbENK5IS63XvDmu2BuD7UvlCTW7oeGxSeHBGZFMa57Io/AMpkAXEPX2SDunbU1J
tnxkgZbemAV972GC8ktE3pi0Nsre6Vi6iXPlTqWTj1SPhUanE/Rr8d6TMuINxzvqKS7TFauLADZK
91awkoU6Fduf2SO+suqX1syxEVjlzB6U3+kJHMXM5Nc4FeuNr7xyh16sqEfM/s3LqPEa+VfE2SLE
aHuGPALl2B46BkNmPAERRMu2mz1Dg3tJO7BqnEXPdMEZ98Rf3i72lugAzxmAHUreHXJydY9zXLE4
IBxm4dJNAM89sDJm3OXgTXaoNYsaPPfIKasiaNjFpQbJeV09zeg5FurBS21O9fhaPF6PDFehcAnY
l5jAlcyg5ggqhcL+W41+yKNkEdow5+1bfuB8xjJPFk8l49TFOPp9R6Ta0y1JXvHI0bIBO3a3lRBM
Kv299LLPuoDMvPig4cwUMOgUjR9q2Uz5kgib8GNUQKsKCdIuzsJjdwOR8yXuwkktgHvnFP86VQvV
LdEHJ8SlcnM/LgrWLIHJI/skyOjRReWkO4850igqly6q38NQr+shTSsaqV2LnTRu5Qp39kZaf4Vi
jj0Qb7VtpffgAFFkj1CKZeFe+wAjY5HJOvi4+qhqNytwBpiTc9pmgfvMze4G2x7rs6QkHOMmnAqL
ja7JC+CjKDX0Zpoqeff8iVy5wD2mlCfZdQS3pZpORq3TKr/DHEkfGC3AOFMJ28BNcUbtF5ite0QP
D07AvS4klR6el7BhKTp9dlk5rEIPbCKTw5LeVXFOFDuozBZnKLBLipwsDubV7E/41BiN7aLFTpwC
NJ0EKTTqouKzSy4y48ZQOWmAR5U1oGKtSZQhx+CYI17aR3ZaMo2042S/CJKEf0/IlFcHV8hE970U
BeNtL/4uXx7hphikZD3uM80BlaTY2GTX44LJ+O+IxNkblfhVKcryf+tB3lYBYuvgmWzuJEN9DrKy
U34eMREVfJNCtCgVJTROaNRqUAfXfdNmvvPuJS8BmfEn4lnQfG8ChOz9D/osvroebo1H7MTvElPT
GYLaq6/8+1TYlJF5LWG8Dvz6pWjAGkRr0NH8sUOBmZfaZp6EvE14kMhvJWFW6eOXvNn0vwpcsZfa
SwFOYdNPSExk+RQw0I3P4wcpj7i95AGdOpEyjxb0aJXCFH/+Y6KtrbHA1mj1oy3KpfUFSnrTHsmK
rO+3s3UgmIqNxEzdrxI+capFa7xTSjByI0CT6Nn61m8RJiTunOiUJIHPOieYWb2HPOtsd4DVRSMV
vqsDlHmMTfqayVnQWqMUI6f640z8GMIHF/t9JGg1gVxdceaxR9Hz0OKoynimHuJ0gsQWFgdU8sNG
pBaktMKTv/EfdEp2JbSQCw8twNcRKKTKyC1y6Jft92nnqw++AFWBsaeuoodJE3Rebo1vW7qQTWZv
crY95gXtuazqeFoyiNTuAwUQaC5DlrPImu/Olq1eS5YPoWhoCR2zELWDn12gNxjXYQYzJ8RhFspe
hZX+J4pLqMZxCUVisjbSiWE3AdufrFsjju3wIWms/NISEJAW9jGYUWfFGXpA6Vfd7bVPvtfzlSCn
a2somiDl0Y/0JvaYvjg01UBlhFpwpywadvqvnnSl8ZXwb5csZ6Dfr32J39Z+Lsn8frM8oWX46hMS
HVavMe2VIhVMUzRCIVbek0kgf+d3QRRvYm8iCNTSiVpPfan/qZrglx9+Tp2/X8N+Rv+ersmrR7Z0
AvQj1FRZNoLg8wkA7dJqK5QgjPAf50rsfgcADX4jr87ULE09YvNQlmtoMaKxFDWuOnaon2u06+IR
caPqIHVcJOX54W15cCgP2wfD/rJX5wolSjo3hIOcI0YGykQIXGHcwWvdGmdxAmz0mqehX8lA2Tgi
SeXHoZDYLxrLZa63OihD2CjPK9yT9bVmuq1G+hYFG6n3MqzXhcbtwHRNrnNC0RTQo+ijJRuqaE3F
oSKLvw3WzC5I5/UpowPxFVTtutGg25Puy4mHQX7l4eh8LGGD0WiKaBhjQTo3/tOsnN59mg0FYSlO
8kyhE4RnBQIZ6JspCI9Yrx8ncs4Spzd7ap2QX8isGMHnlexW23wzQUiLbdvxA5N92ukKffqMmCzE
VDijF0ZrRqS912iDWqaoagJHyhd5WAh7uWUqIJuXprcB2863CXcKXXUWjILa2gFOmDFlinxO+8AS
n6I89DU3SLkeT1h2qcVYRg1nCzZJscVIvflSxFIkvGv+GJBWC8BkIA5gIYiHEYyIQiB6Yix6TGbl
tTskRlRs2+Gq0A0ykMKgOLRpcXzJ+9AmCwtWVZPzYNx7wdcBcx/n39QdGtY/DiYDyZeq6Vgj0onf
ByF5qUmAEG6qYvMzJw2bzVQaoOI587x5dkeFrc2916G6QJHL7d24mmqA1CrNmIAKnyEYTyzJ2VZ6
mey95gAr5f8hZgMtHotECqd8+ZFS6zXlGHMimZnIhx3XumGyQxmM87IMZoTVaKgsFBhm/gQeUmbn
ZWLG5YfDC3yh6o92tPPqrAcCPS37fdplKPJck1TbnaONhgC6+IyvaB8AX9YTTWXiF77DMWiXJac2
Ob287aW2z4i0yufGxx3lTXCBdQHwshn3RS5pOSkmHXX7D5GJa0xkwRVdnDCsjjqL3bF0PQ9RdQs7
n++AeMvo7T7+X+u2+PtNN/sc1HcDrnszf7TP/cNta8nmfKAVy+NpjWNyGdTuoaMrL2tG2W96nOmX
7Ho3py572X49pCaUIyN9N1lrYhtIeytyrMYL96DycV64jfA+amLo/4y3bToMZMtVEZBGF08bRuXh
EAYKX/k8EdFcURmCXq41u8uiDO/C+kl977yLiL2iA9P43jBWLdhfbSf4ALUj99csVeajw0O4OYtE
UX5X8OJEmEGmaRs61NbGGdgYem4HlIab6K/beNCj7UkNvD/nUMR+CP6yTGPfK6fgf9c6r7P+jP3y
Gkx07XssJIxxUeNwMd+vGtvtwd6EjrHsM8oCll42hBl8Jm9O5J3aKm2JTqim8If85US7gE8MbmZK
1FlPBSx3KVWS7WnqWkKFldh8J3dzC0mwFJYwIx8dVicepaQNhTeBizt7NhBq75VGdITB5th26d4A
osFd2Mxt0+QyQUixsB6A8CqEBvcvrPz3JKE8MFRpZn0Op/8C45ErjF81fmkfMkMn4dGQwN+FLk1I
Mdmf0dtxr/nukAogc9nbC9tak5LjHFdyu0gBLhwk7FBnCY01kakahkyS8N0vKmd3PSTWMBotzwDD
gkhWni5G2uJhwYZT/73PcR/6ChE5YzJX4sOtZ8wpTs3dAcF2AI1hmZk27IbxFmmPN6KIzZwvQ8OT
4Vj+07Tl12bHEen+dSoN0cMPjteU4R6oDaJYA9dl24dur7nVhgM+4N8OJlMqLbmJfzzyV5LogyCo
Yz+9ojZfWzYJ0TWP+FVP3uYwBsD8kkMYRmx0dttNGX1okXKYs5koFNKNMSphy5XyE5KbDru/P2QH
h3G8XpeU5nVdGqfhUcpiU8FR74yb+6C35C/Ss6UfdHgpkIFcn63qgDgetA77uXMi6aGmbzRLQ4uf
/CSZdZNKBmAwsjdXkY7d/WFTB/7mBDpao7x1MmhVF2FUNKi+vHsaU26d3dffU5f5S7OiOr4vvuFP
SE2gTs82ZgAH3cKJ736oMar3dReBnuYL342GVWzBJ6wX8LOU4aRMO7sfFZTDPpLGrq4ZA+UoSmdc
/P3JFC7dUPRJvKCRPIYUKtq/FBJQ48NPwNrplAK09BZxeTygzpdR9MLttD4cX60qGCDmn0Vc1nHU
KbBPSsmedGig2twN7MKfWzXahG70rq0Gaw1P7k1FdFm9k8ZHeqhgxwNGuTfYssAApErHRYxt6vxT
UTzSV0iI8oooBwObGlyZalFkyEGXzah1QnG5MMwb0R30ixXfVE86FloJdS1D8tDwZJtEnlg7eYst
Vi6l2rm3B0gW3WNqFrhIY/ECAebVUMZBsKOjfOVWjGwxW0mhSOX3puIf3SM288J7XoNOPd7NFob3
fjqWzQzIHb+Bvid1qotO339m5oOS3r9q+vPUs/OP7161e85Uywy3mP2+qo/yq8/ONdCLDa5VTeIJ
fL3pH+33Lbkr2gDcZGZPF3QR9AiuSqlleV5iDawGq/H336IAS7PyimyyDou3s1E1L32fEZ7nxaWo
pQZANcpIBZCTdgjoiyvn0nGaYOGtW53/exlBT2SbRDfq02s2j1gzOoo9bD0HpIbD/gq/qD9E8hw0
lJ8K8ddLAbBNkMiL67VfQ/s+o93V2yF/mcbj0K2Z4rDCcI3DNWTEhoWEdX/OhZYg8lZH6jSAzqVd
7UP0gj/nMlC0xvjUBZdGY03G4ejF9mj7XLepBkiSDcGeLvCRrVxuZdf2S/JEgs2hij6EY0JhK/J1
y7LO4Pj26MtsjGPcNKQXL1iN3aVK96CGN4Eh29z+vXH95CL75QPDFqItnTo1WyKZ068VhvYzSjBr
H7t242zGa3f8lcviciU8I8U33S3JsEuUYQ6FWJVbYojgYWL6OewBc0eXawA/tiEqU6B5ZeB4Taqu
v72dLcWC4ZyjOjEitAHx/XcdR9U4+Mn+CKTL4iqI3nk5wfRlFAgrY28CS0nTGyQ7vr/uPfQI/+nw
A6zi8OdWRtkFP4loulONBnH1Wpzrx0zZEHce0O8AwfBOESVeMwDHK2Tk2b1O7mzyhNMYeqbC7bWX
QrmunvQPcVcKFtBXdmzmTyDnceSataaBxo/AQEXwnIdr/hb8hrzS6KnaMz1mwlFHAQfcyU1ncnhT
S+Spn2Qj5pvwySqA66F7CpOFATgnbX43VR3/ZCtoZ2P8GOhI7dvO+TfNvLvpQDZBvSlINeaPSBBf
OTwaop7epKSYZ9ikXED3tvff+eedvl3NWdn4wINszPy9VACgIBE8tF3JJOQxZtLcXwJqrZdinHAl
/MT+qTAnOCZqil7gX80G09unshu+DT1P/Ozs3XwZwRmi1yZWBTOzhi55EdOUEgaoUkpaqgeknWli
+5v3jkvzaMTH2nj/6oKG3Rj18JzMLb+JWSKJxnlpM4HS0eWgFG6kT93rIFSdeWEJ3b/CyBDr9418
hIq6TBZ//T3tGN99G8wLgy6UeuQv4Aj/xwb+zqO3y0wVGrO+4Qd5RaxhRIyTHrmbd/wRS1QP6f0U
5DfKIXOH6IwWsXsI5oqZOb39S1zY575ho3+cMjOBHEL3VCSCxyQMin7vEKyUTcUbAxoQkKhWFtix
5XZk9ETkgaUMkEUqSufTFCPcr5bAeT/aoEb2omSpIV1R2+kx9Qxu0MUc/PCVE7rO
`protect end_protected
