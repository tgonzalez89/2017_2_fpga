��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR���[{�T���CK��TC,���:�
&��d!��]9�'D`�"9 S%�aQ�`!�6������V�W�l�a锦E(�\gC�slu�4U5=1�N�m��l�9ў��P���B�@+yg��=�}|֦���ָJ�:	�qv�IV�z�Tz���'=��� @X��JO�f��pc��|Ǹ��ƺ!��oni���D���*��qE���)B�91�-���[Z� 
ǲ�-C�PD�v9G�u���`�%�*[�0%r��ߖ7m���\a�v���Xťfړ�&�f���h���ޒ��<peDn�I�${5��?h-����o!�u uM	�=Eб�����	U���`nڕ�jv H�9_���8���g"����v Yi��׿3��C�ENW1�����MG,�E�EIV
7�&�=��V��]�PR��+y��jr{��	���M̹O�Ǌ�%���#%�̩2#i}j����4[���ά�<����	�I��3�Y�<F��0rf����.?ď�W���Rm[�m;��g������i�qO�ֹ�m/b�3]�e����Â��h*6]�{c������#n���a�>�%Ǖ�^-��KOM�����?pE7���}4�ܥ�Ñ��=�&�wF����_U��u�i-�-�tE���6޼�e��ۯ�M����Kط�B�gy ���\gVK�н���χT�{��I�PB��"625���"��&��9�eA�Lʰ���:i��O4�{�n�8�%��R��	Q;�D[#D�na�Y?���2��֋�@������R�H}dCw�sVRHW�`565]p&��g��&�����Z��nQ;��F3�aA�9"͆0���{�L~��`� ���UXd*�a�V�{M�t��5~Ъ��ϛQ��������;�`�$'�>�����ed��0�ܕ�g#��9F4�ym&��P�R����C��T5Zf��v1ha�ƴ�� ,>#����EOEw�{�<��9f7�����`|��y�6�����F�8�����J��"�&���I�l)|Ze|��/�I�j�f���&|S�8��SV�D;���Q�ϠG6��O�����;�Ǿ����z��0@�Nk\�f�*��G��P궀֖+�Ex)2���L��2���c٬��Ֆ+{���!XC�8�\.%	�O����:���g�g�9=�Y�,.�x�e!�C�)����K�c<��uE�_�S�+��~#_FS�w���҉).�;��d������'�6�h(<G�(�٢��E��2��P��z���
��-L��,���l1�X���x�Y�G�H�^�Ȇ���w��1����Ӝ���Y�-ʶ6�)��=�5��=��7
S]�cQ�4s������(�/�����Ԫ6m4>�pnF���d�怶+�]K�|� ������%25@N�� jQ�*G����VF�MPҳ��R�W(�����aF���ሡ�(�#�ˏʭ]f���C�9f�6�mƾ!t��
���;Nx�����W�:�T*�c4UT/��Rbٞ�{.�Z�\gy�L���|�J����7CxJ���m�F q�z�����zjSF��?�|#��L	KF�A�}�B=J�#;�뺰�zp;섬��n~�f.���5��F(���h�-�1 <�o�����`]Mo�ڋ<�<x�ǢdwPFmǅ��w3MO� K?�-��0��k�Swa��@H]Vʅ�˥����j7U۽�I�N��y���D
*���}�x�8��X��Y��0��;�d���M�1���N\#2QV��:Rz���)�����L�i��#iT�s61(�[��a���_F��BN������!�w�ZQ����R�tX�%��1��2g\�!��c�,��a�5q%}7��Č��wէdo�,K��˱!/z#~�����0̋�i�va���j-���J|�'��ָ�צ!�e9�'uW���q�G���̱���Qq �Rm����խ���F�p�� X�vh0�^�{Ʈ��`����H�{�3�{�x��n��C������O0���/��m*��g�?-|^B�D"J��O�M����W3�� ǊW�%���Ӛ{U��� b-�I71��H|�+����8�m���П�����@C�z)\�9��Y~ �q%Ȗ2�\n�6�~jLFտgXpĶ��?z�=n�)��D_��_��;��w�����z���;��v���h5l`�Qw>��MW�N�o��BI���T�@�ԥR��d��G_����I�%G����op�����������0�xOO��k�4I�+m��q`��<Po�
q���!��8�p���oh\(+@5-y�"�!�R��nFA�3XYi/��,r�� ��d��ǚ�8edk��N�hV��8���5�>w�f<�C�RL�T0JLm���B"���3�Ӆ���ꏤk�#;�w"M�Dp��Ѕ�10�4���Khh�$�z;����F�������H�\e!�`�\FQ��B�@x�Ƞȥ�o�UOFHwZ.��ك�y�������6�eO�'�'��*�9�#�o�qD���JQ���{�2n8Y-��������"�.@�S�l�j��V�j��F�n���@q�����ٶ�JB���u3N��^�#rމY}�,V�nGK�>�o�3�_BȐa�A�t(z��^9o�ݬ:��7z���EL����m���ms�6G�H"n��*QN�~�{��F2΁)��r�BGU	�� �*}�K��"�����v'��m.J�.vW�(;Y7�t�`d@G�ɤ�ʽ�&tA��$]fb��rz�{��ﳂ<�xݱ��T�n��˯�kRs&|�+�~R�^��sO�Xl �,V�4�#�wY��ZG���_�e�Œ�^��Ƕ5�8��Jw8��&�H��8ËʹxY�LO��(�XnU2(1�]&3T�%��YBk��R	�vj�u�	X��l����8D�s�IS�W�4�#�Uꞩ.}�,O�t�]�"#E�U��D\x�����j����fm�[���c�i�<,8�,�y (��KT:e�� aC�'� �����Ah��(�VS̄�I��q�s�E70��-�fV-$	~�2%kGTJ@S�x��\=�~�pV���	+9��J!��}���]G�
o�W�k�{l>D��%��Մ��	x�9���8ZiA��Ć�t�ޔ[���#���7�}�g�-7r�V�.T�U���:B#\��_�4�n�:����t�e����)c��<�!�uv�D�6Ǽ1=�G��&�0�_a����?�2W瞉n�V꘍'�9�,��E�C�Ղc3qY�J�S�A��7N鳀n޳,]rl���% i�J1?,q ��N���"6p�����[j�77�6dִH���L4&9�C�v�%K5�l��Ў7�۳U�P�鮖p��2a�V��}���FC~���i��V��'���n��h���>v�:��z'�����4�KLvFX�� z�??�.��G�a�)�~�ɻ�g�/���Թ��W�ÌGH��klÖ	I��"x���YA��ɸ�Ҩ8��־�IpU�4ž7b ��rGX�̷���Cêۧ�Tެ��)LujF�����W]��,�	�U͊]�KT"�lQ��g�Y��({��IT�;x���ƪ*���'#s n(�Z�0'�<�Nx�@M`��/���wv�3Y��eB�Z���
��~�5�n��X������@w�Ҭ��E�򑮓v���Ȇ̮���Y�i�����:00]6S�����?��3K
o�X�R�%RI��x e��9���A�I,î��yQ��n]�gA d���xJ����Q �<p�|��2ap3�5^��JM�:��Cȵ�/�]~��2��M���z�q���]wY�+^&>ν�������ŀ�?�/¡r�ן�$�'���i�:-���Z�����g����@��V�?1l���ɽu��I~���s��̊Bgb�|����\q��~�9�(N���;����2Ln�^RD�1!r�t3�h1�%�D�7tB��}�m7`P��2��0�0��=�ӌXh;Y����[3�v�̀����S����R����6����^��SXT�?�e,qb��ZĮ&wܽ��=��ƽ��}�G���+B&"����.v~!���B�>�s���/�,Y?�t�ǲ��@�S�2��R>�$��K=J諥-
���mC�6J�p���֤̭hbG�U2=�®�Ձݐ��:}��t��@�̓js�c�;{E�s��b4�	�