-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
kFJSksl7KUdl5lrJXrBVaP4Hm3iP6uPyvUylddkRnGSj+N+3q/qD2VjOhHsgXzTOq9uovDdhNcNO
v/uC63DPXbi5gTDVlO0kJSBsxB/HKK7s4lNSCFZjKGxlAQajCxCWCwMn+KlIs2epzEYGMm4E/wzk
ngSLFAnF3ciw2aHZiCnHcvhPSJr1iAORM4YhbzToEZorYc8MM3yB75hmN9qCha/bmXHtiLYkjesw
5uxRAocmKLm2BJhrqE78FJJWxJj2CUxiYeBVWTXUI5He4CMXIJPUMUfdJOUkc2e8pPj5dCkinStu
uTi3h9ur9l+c8Oyx+g/OAmQFuHOctf8kovr6/A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 23952)
`protect data_block
niWNQpl4CzlzMLr7bLkxCuPuQI6KQ1/EO27w1TQYr9u/xjiOZc+1vMKV/NN29wOsqRPThOE4G+ch
sVnuY7psU6tEMnabvHjl7Zhv+gHP0Ep9zCOOjbLsFNki2kl3D6hMqk89zHszEikYN4ysiYWSPNXa
tV+yKXVTxUoGkgH8T7vR+kr0ISMjTSUTwp+DhpfUeCtgRr4HfP3a/kqyIJAFkthpC9gelJNFoama
vTMhbY5PuO8TmYHEXD0zX8ksWzsWJLPded8hvd3IZ0rNrm17zX0Dzl1BSlAOhmBtWLW8NFFk/J3r
pHbUXDkM0EUZNa51YMIn1vzfZ5MebqgMxHp9PIajtrJYUurrY6b+qCKszIIFffhpUSH6RZISv3W/
3fT5lb8GgaT1sbX3tqkdm4hx5mh20kY/fxJTatNdGmJ3gLLeku5GdPqr9WPv5NDJsjYrFVNHzC1I
LPEuqDKS419PSg2OQFFX/UVFCM6xpwrpuOnr1nHyUshUzATHRyLEgQGYK2Cx71Vfw4eGRhd84hSc
UC06Ylarb/zG+yu4vwJGBaZOccPWJxF2VJn/+sZ45x+EQpAIywGk2qXTzWU6Ijc2VVZxorDIliX+
RggyL6mavP03UsYe5pZ6K8E6WfoS3W7CLZV0AQledzy5wCiFt53+gxB8VTCrctUdpL8jTEE8STLw
hLJdnAx0nnZIEch35FU6VqY62uw+qlhNa4m/zUlCAlLBVBoEx2idIGJofXdX07ZMdFrLLbAGPeaV
X3j0Wl9jSU2djfw0mzLqjD4TBEbE556ExNmrF7FevgvTumId0ZJ/4rSbfhmBgAGlFpPxlVdg9giS
GHDO860883rB6sEyEcPqDx1Ee7bSfhByTJpg/km/W1qsI+Da1+qd2ZwveIK1AN+JqZwn8aZvGHMB
TNQuF080h/Ndxj+f7dsEdEmY8kwci7n88v4FRmlDjMOm8YHK8aMgn6WFi950hUm5hcwXCVsIA7N0
6LnfHSvlMw2VPuJMN0xWE2FwE3MnHmFCHRpSev0YfFpfFqWsW9dcrFDtnjwzJzw95N1deTucdr2j
jktF3cn39m/wrwKsA22TxUjPXpJ4h46juBFR/SSLbKCpnehPgwOASf2t3/plftqEZQvdfCsuF2av
EXydNHha6Mdw8cCjjrk63133GEcUbJJFqy6rMCbLVHG3DXTMpJWNWdWSLCbf5tF944NfN7OZfdVE
FqYQ8WqGqbgI+MdX+DJFAwnNA3s0FD04PbCRQ1dXG0Uc9vPFwyiXr5c8AP2kk1deZM2ndq8bP42T
IOTv0Cr2c2QLl83NO2bYpvwvcfrwhoqJ7O+/RQ4lNKZH9IkUXy74AlJ37at1vjLO3cfJdNJp07a5
Nrm3XPOXgtcKEbK9RQK+LEAT8T9w8fNVVQJsSzlAtBUGbcQy91J6QXztTQiKX+9Au/PRU3dZFEjM
HaapMaqfs1twZtGMGZcTZrN8QSEdfFWHTeUuW8kYAb/5aYFRVhpSyQAK8piRZ5Ej6eYmcVYjzePz
XupUkgpOt48/TCodE5GgCS4alRyBb+uBL/ueQMRUBOXYrP+s2zm+9sSzcP3L+YHv48TPsq4++Scm
kyB7lpT2idzbBCyfR/OO5L3+krE7M7eqXuQMaTE7QSQydmRUxNmdLS995YcESM3Y1xrBYAH12egO
bXPtHglD7KFIFkQmHoJuo2Qf9NutsZOG5sAmTgF/x/CM+Ou6Bt9Jqllm7VVk0tSXvQTB489k6AW5
2MPsOilEBfGktvPALS1lb2QsDyJIXTxwb1mWBEdEoRp8MqctcimIUnxc0bMcZTqGHvEmKrIyJ7Hn
6rsSfBUmywM2N3aELfC3HiTLy6yWtohyf7y94nSjxsp6itzQLRXSFZ5C8fql3YGNubPXXjG62oIZ
egOsTaTEKrEyHwS0+duVhASOow+nSXzFWUfuWioo9IHboblC0/zTBGMKjSRBbIqn6SAiHJzaOmm7
jM/s1+zAt/MjKYvtS1WXckdBTpXR8es8rX50cvLado8bk3qfUoc4CZOSq9+dSK4qebLhTotGc+Zo
N4EywzeAWbRMGdquWTfZzpR5MwNLhmMVVUILhZitfTEXIUNs+2lfKoLMui3RC9z2UnLofAMkziAc
w3S/QZ5QDgFCk6ulVbO2ErfxdPKQmsQryXmKF7+CPsqggDIT5q/pV+H6Ngsy7Zp92ZuPlHXzvHjc
BzOpVjioMqOfqme7TLgvRd/Vny0cAiK7fzssv3i7sV1WkYi+lEqs6dXfwh/rEoP89pvMYCANJlMH
edrtL82aoBAgh+653JCiGCJS4iLbEjW2TFCJygg776A3EWKU+u1G4M88SFYDEeEVwXs8kE3/I0m+
8SdNyzDdIfIUGPf+d80tGWhoDTc4arfFbrbbk+eqz5qayIQIUz9MS4CEIPwcwOSjme1Oy5sI4KEx
1kc03Tp2eHVyjrLNYVoEzxsydrq5yMWVWFsU/BVcRlxz6qo0PTwPYwhctx8XmQed3E5NIc6atq81
RmP4DtcM6hVSDdIy1JrImqMK5FvmBLj9WS6XfNXTvHgBTcv5Y3ec7tOQdmlrnI703aZeKyElgj/7
Q8GKiRDGEw9qlBdmOMKLbhSGvB6Ney9z7KnAn0ZlyRYi792vysQr9pT89Z8puEcinaTz+Ji9jmYn
pZWVuY2OCXoj7TKszpLL5dXcIZF2PEw/5qLDA2tbyxGloq1VHOIei1OIgmjY0/9l4ekIrMzooams
PigAgtUxBNGUPZ+Rfgmk2NuZ4j/Q2LVGBkkxG70GKgbHPWE471cATGfObGogXU07pKhJpje0NvYI
mBjzUwGjwxzG9oZ1AiQZnEFrRA/eaT24oOsps5oKfQoCX9blOLEbXXp6Sw9bmwqW2j1NgvTDJkOO
TUuig8edCjU67K9+dFNl4t9cOc7/cfK+FBFYE1e+YrzhvL7vnvZ4cO6FjX5np0z4iyxGSuY4j9Kx
oetEXlgwxbHgaKdZe8c7lOYp1yWE7DVevXkBj09K3fuyAAzLkiE1K8bhYAgEGfq1rkPNdYNz+u9e
KGHlvKNXtp8D+UWbfTfeinxDDuL2YY06qkQzqWHUNRJ9weaIAuO2DBnyRHXnZ20+uoH+rMG+Fqoj
p/xl1YdV56zu4qOuIdEA9+RSTpJ3TdCQVA3mtPWCbonXNCX4o8p4scK4XZpdCv8y6WUKBIkcC/m/
P28SSJnWM9qpb1WZPVC+AiPjrH0Qt4unTXALqAczDEhd3ix5AggEAmFOAmwN95VyhSzNoYVvKEzH
SQDMoO7+9pquuws6BD1JKYgijnY1nyZizsF3uzEhyTbbsVrPRfc+23E1OZPwGbyQNzxU6b334cdX
ea950gMmLor1ldAiosStheOKS0neHsHdgSj7gMDB04VCQkxmFHmgwG1uq3fGmPpweP3R6qGKnyDc
RN2hYYD+lyNaaN+Hxq9IH+E0ykeVR8p79Cie5IE8FuVQsXP40FickOnQyVbDLNQN+Cil/yTe58eL
FOJsk3bP1ENEsVLGbyNpqSrRKJBIDDO7lugK7RthNwG/2uUuM+/Mtuy8tZy8cv6n3GNup5aL7YNh
oIwz9Kkf0uZmIFvH/KxDUa7RvlJPia1onp5mv9Hc6eNrf+/8NjjbXUPpOk6yvo3HoOKt8I809Jir
IAWZM3ZcOsFYUgFC6/ZPg3IX2ENLJiO339OctRphDVJvgO9iy7+21k1y15tuN31wIt4zfaz6jCms
ECa5zAtjMEEea/rBsylfKkbIgMOYkDnW5N86zgtXlHELYWgoxZJOXWp2+7kHNLEPjRWYkcLW+m/Z
V4ZpQLl+RA19dVIYcEbzd9R3u6VOKvqHO10DS+NTODpt616bZnjyx0V7mtKg9Eygwu2uf18rWDHi
nq9SOXKjwLrF2Xom2OhfgmimLqfSOhmIdGsP1jE0+tJTmHU9M+IFxzbedGSMQtA3CF61Vm2r92yg
G8dv8ZDOYv3kJJoBOHFfLZrCbAUaRtA2JDB52yxm1R3jU5kC19ZuTOmRtXJ69u2uXnaKnEnUopqc
fK7DL3+d3gyyr4RCegMB1T8X9jIdF4gqiwCC7F0LpMPfYjugR5MqGOMYnVjoxKIKMigQ9nAt4IiP
dxuYOsX/roeZEpCNGPAfLTgpefvGPFrUpkXM0QgqzC0X3y4iOI9dbLKjQcOW1Kb7GWd4a+OySQtz
EqyE9ptq+Yos0HznhR7XcohpS0rEQ3dFcxiWRpgp5KFdffN+cVIWb1GvAfsVPn7kWQ/0Y496Ah+k
F19WVWoRax9ZO/n8Zax7wYmRHnxv/qk8tV3Ji1xSo5Po2AEGF+bHrm7wwF3RIZ35cAi7Pd0ISGiU
M7pklDhVBsgjBTPwXh0jAXLq2vzWLM7IWOT8ZfMEW7BUzB4BYQdx5+Ws+ItvdsBt6f/gtYvb1wIV
EJBolcBVpFMO7FYqefe2Vv3quoRvUWb/EZiVj12+eW8d4Gif/6Wbk/d+LuPKvTReq8f4sXTFpmbj
1eZvwVypOotPUjJ/ZnUSsr/qRESkqoN+2c9QETXfIBzW84dEu2M6dyh9H4S0+Gm4zwqhRbq1ZCRG
HfPlb3P1sELmxQpxtbsXLNRDYjh3O61U12nWxNC1UQ2YbUJeaQNB1aY9bZVvVAp0H7nTmYlfwAro
fhByHKSQ9pOvYiY52UE9dpsk/5Cs2BHpBKNDXjjfQdNkAGislOPhWLwXCZGtHv6ZwBocb7angIOn
zPKy4Rwz2KsR4RmwFX/3XcKBEARgX6O6nZ9nF9NDrCBqR8a7WaZkfRGS43RCLklGJi0M3O14ruuR
uPAUUopOIqIzEgStI7EOOtLn2IVhI8Ie0Ef1beX3f9GC4W69h49Uu6i+fKWNP0cHoYrBrrI8kKni
inPJvEfYGLNqJRZnlvUjyh+/m0Pky/rIRGs1zedxFb8kl2eGs0txwp85Qpyegk2EG6a8geM28OAX
jFHqeofP/R4Qq/WQgKuPw3IdSE/IX6PNNoJpclAow5Q2WfYcjqj5mXgtNtfVk6vEm3EdX7CEJcp2
OCm8TnnywAoDRaXHCoH1iAFsnZzIta8R1XzxvJ1DdoRwOHKQ/UJ4aYQPm9+XJ1TsuXr/NJVNlzDC
7exHCRl5Wk9Iee/7xaZKSHUdUJI1zrYM1G5SNWEBdX4EXdAFiKuFqem/EkB4FoHyqgk8nsaJ1253
jiskwrpLahGXmgq8kfGuYoJjWTYKLo8dnScnYhEl3GiRX5vqXtQlYXdHzlVDmVSd4IKMTwk/Vlzs
4JHfS11I5sEiKwL9VRr+uCdrBW/DttvilqrCJ+1N1YZAHSpXkKATxUiph0DvrGHvCK6VHaL3LXZ2
NtR8zjyjBirHBlumD/xtQJjfVHPdxMmduO3lBNa0T9rBI1WAuUlvVW18+Ndai0grpNtgRtRd2bxU
67vPBX+WtKih0h/HwvfeacGmFD8DTOmrO4rKjFZyINVtzNEwNIz4YJoubpWNrb2jwSprSdbnZlQ1
Mo4i5K6SLIb39VXJwUNasQxbM+lt9Q41u61ia6zRcgmcJXuEd2pGZDK75NrAT3MJxdZjJhBhOvp5
6TAl6JYzHA/HAvFjwYi0MO1gsCc3MX7p5BM6M0LEWGbxXh/yO3G+XFow771B2rCPpl2forVZvjfq
EhnOPXXMlQ28LaFOIHkl+RxT9dlNI45K+qmIgpbbR3LL+Q4SmEnUuSACUBZ3WeUPK3qehhphWlvS
r2zvGfw8g8nLsSyZDnYZ3a/1Z3RBXwdPs7b6aathkzijDDsCxNUnxO6a6FlUidqq2ZmNnNnt3MPT
cMaOqG6nIiq5obY+uVIJumu52koUjvPAlDL5BLQov/ZIu/8VCvRsbpaeBiSpFu825QfjE/xtuNj4
E7ttbXJ/Zqo1lTlzP/nvpa6ySeAKminA3FnF4fZrQnwgbufo/FGSL/WrKAUTzlaa/OFTVIEwqEkA
sjL2b/wluN3YonjSQGtQC4dia5P1EtnzRNsyQy0LAra28SNFEp3z5T/bC/savY0YFnVmupBfOPZa
DqDAHoa1D+gNyJ1He+8NI6PZBrOL7a18pYyRTnTTP4p/KUltbeYWkHYnybquY2LFdhpYX0p61z5N
SMdDlxeMZuwRpFClmGCjLejSPEcXn8neKhtltD61m8zDdu/nYAmfhNW7ttN9xT5G7qigQTd5Hw+6
ZvKYgkprz6ajblQ8VtO80vutdPSxBcNhdenXZ2IqjoY1hMap8oN7tXISKZOnalMubC01Q9E3CxWG
4xbdwMt1uJ6ullnyQo1Fo4ECAS5xMRdL7dWDLxmvgQdDPx08uoXW0LhrXMDZwf1EPzk4yjX/sIYC
koKA9J7tfx7iDoKa4Gbm+UBrc0+vLYJ9Lz7EYBEJmaUfjUICB2mz3HEVz4LmKYvK4Kt+WiWqAVVt
DCsO790us5q++31/PJeZo08AYK4yHWnBv6UeiU+JFEIia4ugn12BDi0SrNwrWt7VRUPgdywDLbGV
onj2XiUvO/ymRHv5R3tswOhqpVRudwdncuQUcTJAhAw8D28sAhRmeoe2u2Uc16ErePgZIuWv0CWY
I8pajyNjOdxRoqXyZbJmnTy0rGHVeaTuddsl8/Qykl0Pwy8ZypuMszrkoMI4gksZaN6vOXrFzDLT
a3+uRM7tcR7qdkaMqo4mvHIuVup2HAVy9A5XFMyuYRbiA3XD4KwfH4GkW5pC+wlcb709FgMYBPpY
wGkozVJujxCMBXW60GuBJrPsMlHllAQAi9xDtL9KOFq8Xj4EchRVf5//sdtOG8M9M9IPk1xqM/Ug
srCGPnfjOFBDaxP8kORXS19pLdd1rf3ijM3OV5frgq3RcE37irWAITRpHKpwZBZlUcPiqg3n5O2V
pZIbn+KakTxIbtWWziXuokiXWo5+TAGti9nwSkh11fwEIhyfBE4S2Se2vbfoPLwrdGf4Jzhraadm
To8GMj4IYO++ZvE2BQutwvmfCEdu9VlX0xUVR3f6ysS1Y3kkFVWppwRmiLM1qjS7u6ny62CBEzi3
drxBXO03PGYLCRyqWOfgmxeak1ULSUN3D6/lLiBMQRu/xgI5IZ+dHrbzMcJtaUdd+PI95xBbHPXx
d2fyyp32vSER0kvNO9b1bSGyz669Aq9WktEesUlmk8de/OJjEB9XbrzGvDskJWxH/FJ0ayKOIcmZ
KMUEcqQoBAVgHu4Dz/7oscqgygbzrSOE4Sb/RoycLEFR5PguhkMT1PFYTwrxvfgZSSEDBvg/Orlx
lEQv124XZwMbY5IwsNF2eGgHXGT9ToaMt8pdt4/IlupV46ynENvmFA6usO1Y5NW8fEtgG3oTJA83
5aiyLDbgleJEXtP+qJPhFzXtcyBWwBUshPFktzKRLNHABwQGWUkGxkjaU4kK5PQzvWWDoYHYlxEs
Osl/+U4u77hiR0OOm8glbKZKBF06Ff2S1qsbRRjY13tCG8nHdnm2/YuTxlgMknHzX5HWyc6bPLHf
aDESRR8lGRkyOgEkpQ6+YEjSbcCrvZ7Kk0oagbV8EzvvQshivNM2HMPDbEAPtzgnbkrPO+WR/LPN
Jzo/JbunMo6TNDhxL0nT1wioakQ6OLkf1lIH6v+DdlvzpWJn5P5JKxT0pHqeHyB7AVC6zUlaJ2BR
DteS2uLuh3gVbk1Un79TfEaoSsbzcsI8lUQDZJipsB0gnTP5yIm+8O697+jd7WEAkxf7SA2wG48Y
zCxinE7gD+Jh7uyWJCNqy3Uo/BRt6lVdlbEildUCnrM9ECZF+4DcPOqnjc2HRVrLfzcL4DK1bbrf
sVsq41J8zEu6qbu1OGsSqWHdHc1iHozi1kE5eYfoEhIBa2EqWXDheMXBUyoA7opt1pK3fC++KgXQ
fdRHX+cYovKdxLZfhmdiOOsBBzMaz5xBSh46e7UZxlwF9pVEThtTc7MAZAR3Rtm7qCsNsC1JQUNA
L2qijl75XGxVCtQMv+vgEXUh6zCv6TVKe9tOXvxckJDQspaYio9kD1qTVL4UGoB+nztVRhEkIXoV
LiajfBqLx3bxa/JC+GqhpPKQwrDJA47JSH2p37toBhW4cbgzmkgPuIgih0ED5dv5BkNhApoj80DE
aY8dxBOSAF/2HxOrOtguiO3KbGIx8XToatH4BHBajwuwvbVldYkU8ZWn2zt4L15P3Z71zQzOy0jY
HoTTKVNG5edZWho0Fi1TtLnQvp+xfOdo94lPz3wFrFvRY7XI3XUU0prHVdrh7ykMKaQxUwSpy/w2
PFDKzIzm1hTakzqrL+mFySCb4z1PXHwIBZ83i86EEB3PaG7gYXmWf/Erzoi98SJJ072pKa44nCqZ
wr5aUG3nERpL/+igRl6FUI1l17R8WoCRVrdlIaFOpjurkpnzPVdFTTorQ37lJq3SPLKdWg+LvyJc
6pRCMjSwp3FU9fmtw/Pesx59xcjVFJ0GwYhM4FcfIa1BGjeTiFwDwN5/gZUsaIQucJwkuuHWFhDy
usjDmoLCMflbZ41lmHi4I3k9F2Ib320gLij7bEgicpgUwdLAV+VWwaO/q6ZdNAlY2PteFcU+4ZHF
hKMaTOaqCJm86RsUoae+gp9FU3rPqFjKPta7nH+bIQj6XcpQapso9AzobAOpsrIFvGv7ZqNmv7rp
1xPCBRGW0ndc9DRIq5kHmglNXusfotbeNK6vIp1w8TBfntOOB+2nZJ2W+Yn+DhKLeaYG2nRPHlIf
pBhC1YAIdW4iITK8IMUIUjQxs13Lmv7jWqacaFIhlBhaPrkLKH+vqdIl64fP0xqNP40tH4ayTqha
P7glNANGcrXyj0ehTbU4Idyyn7RuQIZPZeoP/Htz4uGjStG7zOul/iKhiBkuSEaxaBWe9yV/feVw
1qE7aL8l6ShRC2szb45/Dr5fIJ738rrCKmI3qx63/nwBQp0JiliUTinmFiCWMmM4aQzhVhivaYMG
oA2YpcN1p4rpHfUIWmKorIFiCcdh6AoarLT/nqFpxDIT5p0DSIB3aapQrJMk28cD/KDRVurSE49r
ZeXXR/L0vd7xyhgPD2brEsDy5OHE7iIpNj6oTRlbl1kwdznYZbIdmZygx7nnBCVjMSUP/jAMLyb6
E02jzI17KDnlA+qnfkYCJRc7R7Mvqoiq0uJKMXDitTWiOVhleOORblsDeDCbA0KFIT/+4y3zYk93
2u84+nNqkpzXPqHJaJif9aS+qiPTTSvBQxxFM5wNyNCloAqnliPa6P6WulfGts/qjJaQbpDTNtD3
Lcw36YukAKzleNELv8KOCwE3S9PX/FY/kmSQZ2JWVJcwQbZnnK44s+FDjMKmKmdpS7dmk63dCj03
/Im/mUliSZ+F3pzybyEAmLdDYqqkkCOrmEtOB7brJJnj0XMH4BTFyMmKZYio+L0qjkaWZehNhnM1
FBZ7hXtDeP34maTA9oNDL4FBnT2wtJag9rXXrgkdwyngL0njp7fQuh9+3LiQReQElKoPiTud3Ewo
MJEcHXqWfwZpkc1kYpaMOB2Jt5UGO4Tfyvad47fb4dqD80wN8jY2gn32M4e89KxldTKILp+TfHCT
LdDU7UqAeRa7gQ74jKI+ZFhGEifc6Fu2/a19bl155tg/5HdSrHQLu2cuSHmieA6aZLRrP2gpEd5u
ybB+zqzIa4DpW++sV2lRLWAds5YsLkOLOyULh4lSPxGsjCRDFjbUBfMohRjdybz+orMYCu3CiWXd
Y+0ljj+rbHXCebyGXvOueIuHFZhMxs3cmLskA8X3gYbgJxHuxEHSydlotN/uUPctzUQ/B4e/pNTC
4xhtg92FOEYtdEF0ZAgbplJ8Jj/ISOedX4qTwGsun4Va8QZLATLKFXdT4y1lDAzbao77FaoHoe4j
Xg+IiXdDF4ytN5X4r/LVUjwAdihpPHwkC2/z9SjSii76eN1BlUW4NyJ58lOQTz7tiX1Y86kHd51V
EesYxejpltgKkGf9Nk+HfqHFQuIO1BUUXSpgcSAtYotCjWhvFHetNvmCt01n6E7O18w/IVXIgNAZ
AywsBQ83wOWiM0Dv5G4CHjMWj1VihkrpdC6Zy3WW2Qu8BX0avdwS6kGAwHg+nCqF9vGYbKoTaHlt
zGSXpGc3mj+MhKgrd0gJ4MdlNNLNXG2pzYW8KEKDI1P0Uw+iJiQnYL4xhy5pwip2FJiRMNnQidHB
tKFi6dN/MOfgEJcggQtA17wnwaknXuJf4AO/60gASJNLYKM3ocmJ+BodFOkTinYlW9URpACg3zbr
gectFp0stgs0S4dTn8AX4Kym1sf9vqkqC12U7R7sSwD71aCj2Dybo2tZ4jDT3YpzN7epTto+GXYZ
QKIqg2G83GYc//o2V5wcv65vq+7K0xbiIhd5TRur6+rCz0O4jWP0SVZxSosO+966ikxi+WVPyeQC
FGJPKiB/DWXbiFqTLVPRI+HgenjzkjSN8oteTJFSmtfvARrFN/JdpxlgYYfDqa8NuWNzkipOZmBV
mFbY4i8TpiEo3ie18XMGPm5lno9n21W93n97JadSCro6c/cYdK8eiHNTaEZrah5v4hqZg1L8pveB
vO3uBVjeQ0RljYrfqU5JokKD+58D3C7341CkfvdnmqvOv2ewiF8RUFhdahtwF4F+MVgA4FPn6+7H
tT+Y2rLOFKHx1D8lxy9Bj7O+DAE8Dk7CMi01Z5dJCpAuao96tra2OpqAj+bUU9sRF2U+eRV9TvYp
AfX4zGTaehsVSd47E7CvUzu8ZukgUb6gPYoabDCS1nHpUcM/deFvob4UshpSnj6IAk4wgyF6QrYJ
68KfBgbnKGLfuxfh8iOu8wQci5aXL38KxtOj27jbIln20RONN0p4DsSgwSiaRD9oP/Wj6vavOzBY
4zIqhqBwvaIGycG9HRSoIPIo23Z0HiN1HoB91P37cijmGLWfAY/w3t5T020L9tWEiyRh+wFng7BZ
FMGxXCK3F10J3KRuRhIFDjRDiVUvcghAe1EFDzjSXtaStPAh8FCBgq+WQnT6Th/LaMMbtt+WHXyA
iCtgsU4lEshVZdd3fjhpS/rFvf9gP0+sOELin4xOi8V/XXpPQd/zmA1T8OIkICrfRMF2s3I8pmvE
uhA236UzUZLYO24xdUgjT0c5Nwf1ijEnSuCH24IZUrEGaA3UlOw6dTnBDOsxzspHmVXhf3Y6T21E
AVlGQ3yam650pMcX9GtRncuAWfBp72QrLwvJeJY/7IeVJscZUrFcW5P6fNqSfOCRkGpOV+eEqcAI
Th1fXynQJc5uXQ5Sbvu/Nrx3Gs0E0T2DCXhvLnkKTczxouxgP2YovhCVpzGkSAIubCWaEGGlax2Y
VCv+UZe/G/MvW9sdQ2FaX6n3dmexcibt4CrT2dWBpVSPsf5uBBMnzaIoppNR8tIbR1LvzAG8FwuC
UuwAWCbp7c4mWuEIBP/valTs26SLdPMpN5GlKs3q0LX4+z9FrnjzozzbBFR17kNwr8WLMq5JVdrV
SR1XUtMO84OW3Z+qIXUilK9sDbxvlurUMuU9QfoyzNq5y1O/n/OZV+QJUNDcGV8uoHeHIKSF5rVC
G8fHhuYe/xXUP4udVLmacW4PL9M6lsa9IuRKysnLkhJhpxP0Tm/dPNQWaw6SmedIhiM7c5zPeW3D
2ugF+oCQN4mDITa2dTy+WkjvNli6qib1LObBh/9iJikXLA7ehDMMKnEIkIvJu6FGd1s8D3h5AqQi
p2enWYN5iyS4YLsZswyoQijFlk35dz4rseaQVy45M6Es0JrmzMX6P/46Ue5WmsSDVpZ/afgqxJ2A
VU8B1FbHgNVKPseEZhaBaBOZ7YP8S8VHdOEjMsur34JZGzd4/tbACDX6kIGh+iM1wIJcYcaqGlpw
Yu75b+z63yPNOi3xIZSoyioxLdukl7an5IA4PEXsoH3nsOyeq0g6Qs5JVMW4sn/0Oe8PnHL4GwVk
iu6qB3kL4oYsOiUVGagrbIjMSxSzvNv9kfi6PjNgsObCNRUKt9SY4amh5+MxVYdSPaDNQfhB0JIY
qQxAzoVkM+ehDBg/Y6bPkrt4FQc72sooRNWBjccChgAhh13I4j6SkA1tlxreCDAssweRxP2yHcIZ
yRBo41xifkY/wrGNizQxZeckzkOI9oqsuXGuns/FsKEL5nBFQbwauX1ynw9Z6SmkWUroZ+X4/NvG
1jH50EUHmWiJG+gnfqEpq54LYz1qp/dJ9rBss2TQ1HZeJ/vlLBV1pD0RpkwnFInd83gJj+RaBhWu
xqJs5JD5VI42aQqAK8+Re0eWwa3MhAnPVd+v/f3bmOpSDaPRitmg0SSkfXSg9Lm0LyGBFmgXzk7z
0CCgmZTw8tJdVebJfmquOGLOXCCXCIvHmVpjnuRtUH29yVui2e/ZLl2qYoSX4D+fFjjfkJBWHRb/
NXGN3IvKdZEI1zDY1poRANwxeoBNwWqs0gpZD28Q+4EdIX362N+T2kO1vUtdqKuwqt5T+9QSlmqV
ySopiOlfjIpiiA78ZBg/tHjkxat2zoNmFGnXn837RKaSYXcuc6GreWczk+n6YrHXGMOeHMcyZyYf
NM9M5H48EYJU0ekWTl3umJPcRGgKru2Os+7iu7jbkMLscILuMYvQ18j9k7s5QkXwlnfuMdSvr32u
Xl3l0KlVQK+/w6kRc/9BsJSyMZLP8ZyTcBAnLUg0I4DCGrf1bWslXIXfsX169wH0RYiTaNE/r19h
/uNN5SvtuYJwISDty9qkvr7AqEFgYKf/cOIhMHXLYLNbAcwkhMR6B0oRsmg3TNmsEPbv4Qxl1qH8
3RYMWPouB1fA8Mf06FJHYWjp75+6OUCFZSORWnuJKwjtKY+lUP4TwpqwCtHSR/VAHc2gnAeQy94H
n/CM09KPILoPHJiVXZaE7U2cRrE4SzdIrfIW/ubrqY+gsueJg0YshZO15BXmiXC/ImO/eBDy/Buu
CrZvR14Kw0LFQ0wYB0NVwsrh81QHrbgGuZHVrbTdFUyfNXeDPu7NL7NEoD1RgKncxwy2vxrCETx3
UZs3AisLLzIFVWaFTcR9RPoYH5BklhPb9xLK1fw9cvvk8zj7xPX4tceO2KqIGBcgg7BBHxaenLmt
E2hAcO4b+OUE7FPtYPLc/gzvIEnk8eVdWXEVr7A6JFxXCIqHWEgKRjSVVg0uX8Lr3H7Vxy34aHev
+RG4IcwTCTOmXLgubxlowZHFw8yPaBi2o1h9R7rTn0I4pS3dC5v+GMLP6hf+hrJr1tMJvyRZMO/9
xw7cP1ba4SqgLwzORWdCamlwHDnsM1HcFwYhsi0HqIR+ThiWCsU4k3z+xXSaDeytz7h8gFBhGwkO
5txaT2d+kc6GYQ8zFldNQf6A5IVOjEW/x6AaSfzRrthlI7NvsJh5NFWU9eDzN1J3l6b0eYcgnukm
4LxCfqlImXAUR11FYaLYTAqnc+oIC3Zv4zPsDqYB+SL30Vp8z7ygcDgn5emympkKXf7onwZrPLoB
tmEheFlxH3rP6k3RBmIvfaNEn4rBf2CyzVSurmR1bjTIl1H3ll94lkdIP/nSyX6XFc1V803GcX0B
EaEc0VlqhewfrN7zo7lYVn6ArVGykr3WJ5FmDRxT3E8iwjLHQxH6IFDk2uEA4HjnkcH9YMTUKV3D
wA+AKOQJYDJLdtsQ+7XWpcRooPojK/tktANrnuqKrBO2Dd0luMBtnSuDvdPBepoH/x5tlpaSJ+lJ
6F5KMX0xpBdAAuvc9XQRjpyvKhCMInb1a59rdwnxhA7f9IZzrcjvbRD5ot/0BFj9oGO66BsmD+G6
lTCHnksEyp497xkgn8IQmQGEVJasr5RP8NnrIDRI4Rt93X31CGm/TibrSW9s0rEy2takO/orC00J
o4TsPbJBPrt9kjg+P8HnhZukTbqpdEkYuxTDuRdx4ZYWadFtH7Vje3lx95s01YTem03CCAXJl+E0
MNXR9InnGX1bi56Bf2xaq6OxtO/pHMwcVEhaDWmzkm/WrxMTb9ervA78M8SeVgKLMkXz31AeJ/r2
PYWQS4tIU0Uyr0taHichVl1HNwCgoGbTw5TtXZbLqr/KKgAgR8qw/incslbjkU3UapqYK4H7BnrO
3iHye8R0wuTw2oWNz1LjqlumBzNooInA+w14d7IngBTvEZ01Ej75pt6EInl7Yv+VmX2QEMxdSZ4w
h4FDl2dEqUgmI7EXlGMRR9ykDRPUhtcYsZHyPZopxXP0WrNlvPrvNbjidecH1UokCKp6+1U4W+jP
q01N/1vX01AXfRXOuMXt/HJBc7on51xVWCsI/hhH7M1cQs5nOCfJ4g4Kl7bVxCP/qbqoyHVCOP10
k5b1ZFfFUX/Nuze3FClmhzCXpJiXth8WG9mVmYD+JDaM/3BkVsD5yO7Y/ZHHR7en1E2nZrY9cAbc
Wj6FIWoyrGpayt3ZIMz/a22auhvx0VIKW5zHXpaG6D0oDmKZLlox20O7DKYRAcUm16F5ob4KZ3he
sgoU8sM6uQ7URF+0hP+0vbA1NGKxyitqkCdijZBpVfDuD8XEjj3pxPqc8ggjlO9rpQyUTO6EMPJl
BAL7XfQD075l7VIyJEwW0+PqzGh0TIgf0WIGgyw8Z2SUJzlfkF5zcs4qvE/gFB11RNYPFliil64s
e+FVmhBKAWitRyHHvbeJedFOjpTQGArSom/VX1Kw7y/C6UFN3gi9b/GQaNXLz4OoZXE1ZwAQ/hlj
EhsXhdPI6wmwg8zWy5Uc5TcGTgF+K+GYHqgtYqHPqN6bCtnylKRATJI/LPmsma8PGNlkC9LQ9DQG
+p+G7uhHK1Oxgui8ztVqaU2Rsp6NrY9Qc23CgfThYx5pk8XQNBlAdUB1A+2XZR90FhqQrfddPF1y
eAW8qfK4nvI/phWSusWqyzHzAuKuRfN2cl4ee3GP9+tfi5VUGXfOiBphAyH27sqOnS/5nww2ZW9I
dyQGr6oc/dMNTHbgF452J8zO8ORFNOlBRcrz50BNhjqcLRTcRxoDkt76nA4TqDdHuv8yg8+I9SX0
Qzor1UjdxjlJoD7Wi5cRbRNUt9dkvxjkpHE8KImpbzHrbtNz4Yfy1V/DMLkPdvt2LHKted8kt/KN
mdN9DeiatQkZnARLTu6kXYKXI1bItSaOX+C8DUh847eFzG81bRPy/XDw7y6F4ywPZdEM/USyObjZ
QgjwhDlG5+xrXHSSvFhl30FL0I7kl2An1TC9TZILIKZZuQgrmU7OguXCUcS9BM3VvHK4oi5JG6ak
GEt5jfqonqi4LSS8FRn14VAz+6EJKKiiXuMCbO8a61FZC7Pizdd4o1FvTHh6uozXiODF29L5Qqqx
KhpjWVQzp5ByaiF2GBNVLNITzgORSJRZtoUfUBsunx1gW7sWsK4b/j+5hjgz3oyG4RsAP3Mb+4Oc
913C+j58mrjtMobELawLWZZoZH2vrSNJnsuDHat0iBaPDQDO1ZfIH2V9S/1kXXCvlQH/XXaurhJd
bmLTsG2zVNViKi53as4ahVsst66ys8FS5H8lvNwUHYXmJeQV52o4l5XAD8Q/Hs0pyZVVbktznny9
sJTkMvchzBEiIfO8ouyu3A/5NFQaFw+O3k+0p/cyRF9gDmLFBASjbGzsdIWQgazWSn1bbjstJPBV
7knMpy1/UavDfD3StLRF5HS7PTEkXrQ9cF7K2p10VAVGUjizh5pIWJ9B2vb7QcortvFKEDP5LoPG
sd+p1lX5ZI89NbUCpZWoyWotcGacsL24+2AjhdNODd+YdePluU5giUtJIlKksphlBo41JBRHTOZK
o/pISuGT8xk+kOP+vpolNq1ijEN2XS5IivA+APtcQT+ZlVYI5aahl06/1p+ftCsKz4/EUg+1tK7n
FUxWDzRw1Q33PhamfH07U/23F03sirRKPNX8LEDpOLwlkTJ8Ubkcfcyf8uUsRG+DPNkJYhBH0+Pe
8jUFs9E4Ltwq1g7VgRDv/egcSpgbPCCgR7JulGsF6lGWLNUce3pE42F8kdXRGoBGNbJ4fgw+ONMs
0W7Uuy3clU5S+aRJaCFqr28LOC0twkPCDSOfMSLx1GNcfCWeGIXx2gdQAzO6PQE8r7HZ2m0BF59t
gr+iNM9PELJPIhPXpNOi/PNL7O568KsIglaZOdd6PbVqxjF8cpfcbDJKxDNQdSakiQnvq4TuCqy4
57Fo72xgtyQr9rDkGJCSOAqIYD75Rjqe13Xm/qoSD9N6Cw1Pm2ADzXuRw4gHCxKPqdAVBms7hcdP
MLRgpdaMLrCo8AWC5cq5Q/PVK/9sh9wI25vPTJIlKfYHKusQ97mEDqlN9K17e1r4BCt2oiv/4B7o
OJv39+Ou8aqnG838czPGe71wk2plz9Nm2SIBhN0vyUCDIJ26ki/9zcTU1bI4Q3ryvKWUE0nNAyag
I40fYt16NWke8FXJCu51H5x2W8o3G6+Y4m2dUJDZoCYbtnA+0KfOemGHu+zKlALyVJDh7YnMOrv6
bCS0Ehq8swhitB+n0bMET2GwoflSSQ4vyYzFelVfeS0fEqiwQu9Rcshsl9/FPHJAPBmAIa2PTLP7
oW2QpNAlBYUBJQz+56YeUkOYFSQa77z5y7dSMQgJTFHlH5+xmy0F0aU9ZInzPj49iuXWeDiWILJa
NoAfy5OPMjZSdzyNe1DpQTHfoWy1B2a+IBrWhZ/wgx+kTouefBkrhAMiJP+cI+Mr5C8Cxta1j2zQ
WdTmo4Y8MEPAptpuD1u1G3ess7lcsbElpuK10kaSZE76qCQ6j1MG5FfvAFQXEPROHhoSyv0Cccfo
oBBggcLZAiCJ2ZmfJQaXw+2VT4LH3oVgZ68n7uAxAMM4ir1dObcS3enfKq0V2yKywfI3Lab4YYBE
liZNxn5wWT56AZWhcearopCEiCSx2IXOmz5Vy93Jb/BbK0dfG0K6SE+wyL7mwRL6+C/abYqW3vBA
izOZwsnxj5gPBOc5dyQaA6utW43AUFEPF9N2YfU3nw21J/QU++jkOS2hlZWg2g5KBii8DIAJnB8x
HglD8eo1p1D2u8pt8yOw/oYhe/zT1NBc+uMjRie5gQpS8pzVo8KoTY8wimNABv3s6T8iGQKeo4b/
1HSdPaEZMvOYkjBxDh49cDtECzgsELbm0IKKLanvs8I3UoTgYLXCz4rGR5xhOQZ+hhcPIRDzVFrO
1QsstRBkwsUYhDc+60+a4Aa146ODdZ95RH9MFKQSfMx1Q3GKU5+rdMyXUfYdX2O/eJf3PR8FONeu
jQ2qioDk6zQuq8P+d9ifEderkVvzuOmYWio40Mv9VhMmlh/rTyX7kI5+rIyhRXGXfanwi25e7iND
aVsKhceJphS4g93+86vDDIOOkvMx/OeUbX+dXKZ/UsaXeE9oQID6v7PS5JhNmyx7p3cOnJyAza8g
/XMRg8j26IoISePvs14jyR8aFA+eO238nvabEE0XQu7K3nbv0/g5XPhmtoxoI+5RGxJLwQLD8bRk
xG0u+cJv/P2Bjnm82AaDL13GqO62L1R1nRx9PsNu6SnDS0eMYz8pSQ6//xgGFOQs4uW2AVixe51Y
6zucrm1g3lw5XQiacCPLWP4o+AT4CrUh0MWwiJeZL9zxgZWSfhK5UJcrqwJnw2OVSMWmuTC5BJVc
aKb+xRqVX/WnxRj1boWxaTlCFz0X//1aLWbPk+78FRyv0/yyMuDP1SEPpqR5lgb+OUDsnfZ69191
r2y0EzN13T0RXI+IPYIA1dNJgCP6oPt2O7F5LgnhvuqIHpJXyI2hV/GGRVi1axdpBox8GeDuxvKz
/ru+rfphQyh+HVpYjuXtE6vfbiPfWlLwA1+5ggMVPPZh4urb4EKmWnnN1wZY1F2yHI41SkieoahG
+rTvrS5IYF8sFrFSop9A2EviLpSM1nfD/Z/nCjX8sqe60SMisf0qblrx017Db5BaSLiK+17oXHKS
JeRfpELWsAxTn6twrxo9ZNsqffZVcj1Y6cA2lxnBvRBZb0yK8QjdZIQNt5e0P/ZDf3B6KmjVSq5m
eCnWUKUQ93B63jEuR4n+cdpdUULspC2If0GIqNh4DTe+ZB8a42paws9ObARTLrcAxfceLjxSw0em
paGLR2w56GGPPW9+cJKx6Ru3qHjfut+dvNyqzCoHNUyGlGEIU8Vb2Yh3nHrAcC6UBIfzTEkovSP/
g3wklvmnymHVc6lvob2tUlE28Ed0kZJpzKGU/YHV5Du6F/2WN0QhP93vzwhoqyJtTqyRW/M/cTjq
+VMCrIsBmnzpRGwRtZAvTEZA9d6/IHgSKO87X4aIeBvPe2j9sLI8pjVlDp93ki8HzM4XY5FRTpBf
o01XDznXH/ZW4NmiXLprRrVV0reqIeXqfKmLPmYHyUeMlyYm4Awgy96JmKuFVgJXSYOLcyf8tVCg
1rdCXweP/X3hUZB/n/hDPocFjDyqOz58IXp8AS1l56hVBJIcCIrDRnrkBxY+3gnFYDGE1+f8161F
6poaJPOSZOfkEkDnnPWnP2XgYhtt651vONBeC89tYjMVJqKrsPKQ1XljcZdxguMRPKs8vP366TU4
em460z0miO+sHi8GMP3pKPPL/qluKaICfOB4QDXHmlcB0xR9cvDwMeMVQLPv8IWLZMqMOQez0rKf
Ffywd6ICR/6RxdCF3zm21l85jyd4oWoZjM8XgCCWgG5iWV0W7ZbVVDVcsArVXhRxU9SEIpPn8CLJ
PHEs7Jf5oQEcvEKbTWi1bg7De6B9VKTCnEmzW3qZCvEX9CQVsSdrADfBQgWjgDC/O3J/AA2pTQlb
LVAYeF8lNtWLpo/0TaInpw/q74yuFac1mNFgRPDJmwfYzSpc5oNP1i7WDO+mEwXmbFfvoOxOeCJp
6M6/tn4ueT9CLRUcOiOS2aw4CcwV9TfZ97FPXk3yAFTtaQTsY6LsJqv9Co6P6MLqwokLAfhb8Ebp
Va3+2Q2cpAFjD50i0IXTOPD/x6PDO8fASPpShrnUY5nmvndlEqPJASfp+MDzIIMAu8eecn18LNKR
7FGto7IXr3EdBgXveKobqZBU9/aKWTe6Vp8OUEb3x6Mkpuyfl2M6XKoBKHSVm4s6ZRHWdck+K6OR
5IYiRVSdOnsMMcZjS5OTNv6txahVistmAlLhr7bUvMo1L7WeN7AL2SFErPt+Pv9DpURNuXJDJKrB
MmN5Q438b+0UA7WHLA4yxJ0bz0Fl2BXgXKlZzu405h6ZVi3Ep6xOOYW00IoxL7ve/eJTPlL/MZas
MwHb7AiDDE6hPt8kqy+nD5WKAgzg9LYjEmPSVWbiBm3SZShd6QSL3Qld9T4uzZxMFSUzDMqsG4vH
8bdG1rktnsHtAtzrFCoJoYFyhD4xm1aVfMNHIzVSln6J4RK/Ze4JytyYwX8GKBdiRjWjLwZFuWEY
gL09x9fcs2M7tguvbOeylK51TqVkcHb6zWpYXInehYtko3YGq0ohlChlxkepEHtDFUbHxoaXHe9e
5f+qAq2xxfwD1vScT+zYGn8N61cznslYwmZ/3Slq6lXFIQuj9D8pbOyR670QdP5FpXQJGcgH/ku0
gYPN/EAV7XKCDslo9+BRnTK6z0drwc4VTGGlWJYWqK/ZoViLOukT9mzFux+Gco0Q2N7pF2puK6qB
idWslmfk3eg0ewXYQYRcSG7lJBZDQ4K0WNP5EI+PD9c5Aju9FtAPlMzQ2MnpLVGSVJgNW/ybcwaJ
SJZ6107Z9z1Zgkkoxm1VdYcmjKC5rXbWjvOOU5LIL+P/x705GEppj4ClcfC9sIALwBlEkqBxxGS9
DhGKqEo1v91J9Sc+V/fY3DYSav0HlN8DqlehwoE6uFToFrUOlveIsQuVsHZAzLq/MFNbPgd+WJZ5
/kUboEsQefPISDjfacfJNFM5R25Go+15qJvSZBBC56idPg/CiGF0nVbMUttW8dzJkOvCEcmH7+re
4XlBtbb7+jJ8/7XFTUsu5+47hsOOx1kGW8QZafZswYoeJj22UBtCptU4nCqk/t75rBaqpUHfcEBy
+/tTIhJL4isa/Ff2+6dYT+zpQnhTEK0JDfAF0sWcOqvDf9HFu27FV1YNYvK54IFwuSu1MAq3lTWp
KrjkHUHQFPkbT75DPDjMyaRJ5HUySN5gLgJ9qONbZOBFzk5GXZ/b0HmOWAFyAkJyq8wKLgMC7irG
RTsf5v5ayJ6PqrdrDGYM66KRPCNat4oNO9aQPzAiUADPQEOO0g2SvjBWHjgEWojXXUjKI3pvZpWA
v/1O4L0k60LbP4BAf2gOq3WvEzLIGp6aVpa6WepKebhCt7BF3MxkT8S/zKIGYq6HcY+kyw4ilGYA
AgxvP5fih12mb4KAvCypVQwDZ3dyI0tGFoPLCzjpPlRPisfof25n8WkHlysnHpBo90FwERVMAqIE
rVCd6y5HfBtl6WjrdRvgOJS6LMIUM2Der1NDZjEvhKTwclqMFljXXbYMbGrA7aPUndpXPYlMNo/4
0+bjvTi3NNHkExM72RGMBtVt8NK6BdXIk8oHy8Jh29VROpXHWc2ilMwZOSXaEvFmwBEeYQRjTBgh
6YpIOfgGgqkBjnswRyC0N1VaSgIijOQmQ1saopLqs3/nZ1sgQgtYCcIpm+lnc+kXFuI5Z74X0Vpu
7wRVebdVuOj/7f/+XjDPJhFWlisq9z1nasJrlerfkW7kK3pP2UUAC+VPgPHVxx+fIUpgdHnEibTz
dWhb9L48vVwS5Jmn162EpXRBjbod/A50nocnKaSvm9CeZ35tuP+GZbGsGjdB50rYaUQFu7TT0F06
lackod4aFQ5j4mXkdotUi5Vlev1GQBJ3ltwIbuzw6sFYwG9JKM0yvVGZ7LtzeTWYchM6I5icZSiE
DvFRQXmtJizB5EHAfn+wosjz9DTZAKl7xes7KjdIVPF4P1u5yzYD1B+yd5ZKQGuXhLnQTgTNd3Nm
i4IwwawdKDIVw+lJMdpWbYSKD/5R2jke64ml5pEcTVRbAPEers/JlVbFq+58gR6ftYfVAN7OEIMH
DZoj0spqHpzxFqJbVTUFFacPvJHth6WPOpAHD6hX2xwQt/osQljOvGvIpsgvQxvQmz9X+770RIVw
xCPlQTul9a8g7Lxq0SaceSiXLnREMEY8d+LYW8xPzw+X/DUGo04XzLwkLEeyvmkeUDtUWVOX4vSM
I45TfJ7l1EDY3+dYVMDs9ClTiwj3YrwsIRaC/ZKtft/UVA+y/Fncafmom3BnOZOWkYxOVIzisvf/
42ngZnURcGhIjhOtReHlYeO3HK1rUklasBJ2n1E8yHR7mUqGl6ZsD4nAJLz05r5R+bbW/J7im0OO
xfeR4hHmT2D5kqksuU5+NMrH26X+GXp+PfQwoc7Tx07asaf2jEGPmBlPXxmVQKWkQdJd/8tXuWk3
jxhY6z/Wm/EOUCVwxQqNjBe/6f/s2DjjIUDEmGc7Qa4Tl4kxb2fG6+6/uelW2ciDKobPIkbxtq0M
FmNHoaeUAo7hK2BfVEMMvTiZFyy0UaOcbRyG/ffnIVq5St+Pfj4Yrol8NCug49P8paH4FQYhXVsY
L88cf+jZObCCA70HAP/rVmt+olVzS3QZz6YYyfMyZIfpVuJ4ohJ1JQKnoMpkmy4QSdV5+7mdfYVY
zZb+LMipiXxm73E5wHOcPKt4pbh3UlncWYWnoCFYiVm4Y1JXztnraxttCBpFMapAu0nx3UNndhfa
cJ7hmN6E3ccv5J4cQ9jjgWong1BV0WeyqwC4GBqTAI/ppLdSVtziuT0WJLB4CQ0VVkXODF/EGa0Y
I1P9V7s2od0bgfbWkVn03hgl/ObG07lMnYolbb8CiXnTQb1ZbphmkYh5Zfc3AtDHBJsboMRkISdB
BJcOJvKFCoGKzI9PzQepJtNcn7FsO4q6eXgyyaLTlON6mjj8vQCpGGmPLdShnU5DJnD25KxK53GI
aI/eK4d99uWc0I0IV4ucOzeOertm3jDeVKrPaqo17yOf6utZmkxKw1RtA8064OFAcY9BwVEv68xX
icjwgWzFQp22rzIDM3MaWG16AShqF+0DfuhXZ+RJZ+ImtUlqLMXYJMM4B0f5MrykULPd4UbV6Noj
Uq3xqfQD8b0dKNJXWHZz1UG4rXhpwjDG0aaLu0nrHkdlOQiX0GipW2k0QZ7ZJSXs7q5JU79fU+HS
6ACFVKfOGXrLhLA/Nxb9JeLKbMoL0DUyF9xhYxT9F5hQinpfVdfVvTUcsjlLk3twF4o/OqeTLHZT
/A/vB6ELWLOeBkE9Xc5EvVSpDV692jTQfvrQeAasfvGICNrnBWwxhQ+xS7mFGf8BlPsEctBLzzu4
Y4h1MUNy8dZEJPO4kNQlDk8+P93t/jJlXe0Kqec1FRC/x++c6kYufyR3fttWcvkKKW05slX/5L6g
GGR3m2jGO66dyLDXfU6Mw1TIGJ/7EfXyYMZthjh+ghNbjK3nBeFJKMGYktu8OP5YQp3gZplYeNSB
Fsv9BZSCxU/pBd4x9ym7vtsjdmHvltRvi+bZq1jR6Me4NsT4axA7f+AR7M63JSShA9bsTCFrb5dc
Z5oOu9gfEPrEKQgZRf9X1snmHOsL6kvs9ffdiJDFlnWMz2a/MU76SaQXmkD+hu/cJHpjMs2/mLaN
i962hc9JA39kc1BHz4q2mkL99cgIAhf+iOKXcdlVhO+MQkd8C5LbmNu1LnZd0Jn03Dru396nOsN9
rDqdgr7wCcsqvf0gtT7fk4iAL++UOv5Wt6PIitNEBt4mXmgvhy8rcoNBnFghRUwcPTrknzs8vPCi
XXbwgdFBFMn9QXKfHIlDfDZ736WVVUX0pc7rDb6TUf2g59VUYrkpxM8l7JsOUUWZuC3Ni8ggk6z1
lUJXTIZkwVm3NpFbimoT6qPxSoWN9VZ5OndS2Eep2113sgzMBSFmgg1ksDrP4jljMtpS7HMjU6ga
Y9+y0gC3x4qcJ6q43CeZZJHLzLXFaGUvpj4Q8/ZmETLu6IgpPUIYjNbtY/724g2nviO+e78GvNq4
ZHX0cbhrzHcjg3ZG5zshj2MZMbHnvS4rV4dWrlt408zMWVQBcrsklO61OG9x2BZbIo4I4DbBlC/1
T0dyTROCwUT6HRc/7H39G/OOxkYOAUJFDB3oHRocCk1/umw1+dPI08Ai9Ux1umn8V9DRP5WgWBwx
U96tvZNKH4e8EfmBhY02YAKkgsjnE6DMi31oA4j2rj1M3OxrB/3FH61a5lnQCS6+zvKp+TILA5Cf
c9Mr8K0noASj9vZFD7H26KmhofM8kKRwsmmEmJUNVMwU7+iu+HKDUcNtYUhQyJwKMWCELFtI0pxb
atyF2WGeR3rzFhceu4Jx7e6shR4hCXi6JPadtrPG6A+iFcPMf9TVRRi0/t01GE7VSog5VD7hF31o
/hFz6EAdc/0rTIMt0z/rsp1GgrYtBWf3Jf2C+mSWVu1EAg5EKkkRm8XCBEgxvTEfTRcuk4QDJu/2
zFsMx23gtpsZrxim05a3N0SWdisfzETW3waoT+9fRgrAYjzU0jE/qy7y2snSe+/8cIkzg5vXVLkF
0JQLZcBrtTV1Wxduuaz/xBa0rOh83+XmT2p0VGlzgIreXocLtTH63B+0Z2pGoFKLeqDB2ItxbcYm
lXqqvd8L71F12eDHjDfLIu14DuvS6tMg7pKlPSAW/ZfHdH5+waxmgIEoE8p7vXYM5l0u2L5lGKiU
destkUEIiYm+aY1xQLdu3QVjvIWl7FlxHpLPjsuT+00QyyBF9jivPyqydwx3FVXO5FIhDPLMzgfq
stjJSWgQru7ggWuMgYIgG0pL1a1N9iQ/NIMWkAWeeArFMnfG7PVXdOuI7/0a+4M/nSSqwZS0vToz
qZ2sHqtnpF3EH6C1/GGp+yCA7Rp+bofCZWAcuzRSJquMwHSGRVaB2200dLmlVxxK5Zdsc6haThRf
tMD7v0WfaHMOSsL6D7YL/3b8Io0IeblY1WEd8plXdOE2I6CJCDh7jvXOPjuKSVO7atqZvqexPcX3
vRBu4HY7H1KTjnREnaN3CYOpcRJ6x5wdMmteYgVkJlaBy0faVl6pDEx5s7Ap/HWpg5vWV/KU9WIy
4ewHwg/TwbxTrCflxIGSHlSZCMphn/0CvUJy3fXNbH67UMEK/aL3oWR1OBDbaMOBhjOlBUQ3OWgH
hdQmTWq6eT5RHDZ/gkirleYMBqeliRwIZ9QMKC41KuiUz9rjAGBqOa79qAYofZf2WCxwbnb0iVqw
2sh1CclKmXH652UWFRwch2u4NUWGQhRCY5xtWgbEWmv2iw3y5xBmcegTCtz0KsRtT1R/DFMGdS4f
VHaLgAsAISGqKW0DF42gE5bdFfJ0Cj1h+zTykNhqIBhyjNLJzCgIibEaS7DBKpx/dgeEbUitszxj
qqoYyB4srmoqcc6sx0Hww2SfWeN+/L2iRXb5UfLECtNzRzUZjrVJZtXXNj7aKlYvsfnbGt3kr5tP
JjWEl6dj2QlPk2QtCQAHwCBxpLyNSFGOH/EuDCDOwParUKEmhDAZrA5h27pAcLFUJLVVpzHMo5RT
HXlWLIifrJV48Aaf6WK8KYY/TPoJXUjt0OYWQcZmO7xZB0dQ52qXyF44L11J5wbLW02yGEL8uDXL
0fgwoUX3tuWUducuURwGDBOk1/E6JwJvB68HU9EpBPyoYwpkVyV2vPnvbIGXCRYtKYSJn/xZ+WNa
l4gZgHk4fwDqM7EHZYQvmA+BnDyR/Q7OJ51X/bhsyNnkazgiiBy+SBDw5oDiBT1ucXicebqrxNuh
DBEZxrJMoSP4jPDtekqA8E8BKK5m02LISdLy5elBjmYO40UgtF6RRFT3hEdtV79SrsjcWWmtJ97y
1evHQPvIXI1asIkGFZ2gzl+KYI+/8iD3A6BhNDgsG7skcx8YKTbAjc+4EWhOchTX62UXLcXjahqL
a57xLO7VAh/cu87w8yKrzoNbm+/mjscdd/E2em52JFyY40kw4dEJR110nuDf/r7TyUQ1mL9F9RIT
ssUS5+r0TLgTR+Gv8FVYQ1oAqdl4hFaIAQ3hsRnAo2bi/sqznp5pTmtDLW+yRn88wjz76M9dJV5X
hU7ErIvnhRr7aAR4k9FncIJwUsvrPflE0GBtvbvvnl2sGPYJLtPUYOQ1ZQenPkeAaQ/aT3xH20ge
fcW4U8HuFLuo2Cu1G2eF7CpdKg5ZhSkbxVhUMreLpnPu7B4OMzbqtWuJlYzwutTYkioP8IrspWY5
vk4gTSrvjd8D4DUtwNsKbKcvJslrmgLo5oKuXXFMYsxtvP8+tSQ76ICTO/ZD6ih40vMD0UCm7W2m
00EOqIRKwz0Vb0N6jKUxYteMQxKjuHyrobRYtqkQrYWHt6atxI9Ay0mexFd4Qwgk6xH6SycmmQk5
rXKF13nk1LwMi/xCVd7Pb0I4B97PYQD7ugaXkwrGshprNEvXRJN9V1tp3qw7fXlJ1ZShblUsyNTE
ve7RuLc04brDw8FdYaG8CijvsFZfggytJTHwUw19P0h2b0VeUHyM6VoLFUGpIRCpCioMLRqtMfjF
X9K6siO97soqj3aIip5RViN6JCB/PukZFVxpWc//xRZ4LUPmsw5lTiqQ3tSzz6JiAL3enVj6XTpu
FRdZOdE6mr0kHlDpkAw/fUeUXz53mqQT397zh3vEGdGO/gnCAz9cI1nKyssDWtyS8NixhDEIuPlu
YPoslLK84De+zt2decjONEcTP0JfPfrhGXLjaBYVVK/Uq77eofBI9tVIeYtPLF8xDTcIz1wALCCv
S4JTxwArcRQqxxlrBZtPlnPSKu00yNUJRZYLd3wxZpW718OjFneYRLt/39lZhWrbCZiAPljP7xz/
1oNpRSrHjmzCnBmm3hNWClPLlCJ+VRlMgBxMJionLGDkHJDUj3O21PGhIIYjCv0MQ0saBB2SqjgG
Rc8cB2zZMVvnZgcF13JtvfzyQ/91Xm7tJZZGt/JOEgBcht6zoCEMX8wysMoCAVOPW15jvgb9a4oV
tdKMuiqtOLWzaLJN5WRDRGi/90Poq56PpGFi66fRD/wiaY6Sx1qRk8c9w40LzSgfrjqgOvIo5yQe
dXethtlJjWQrTFailt4ioUaLPvKleh5m+xBOg2b7YSJ+yRIyCri9CQbBcmDPCMfnTiQj6U/racQO
b8TOxpqfBs1QpuVFf2i4i4MPZGa1DVpV4ws4nnhLKCg9KTwuTIRB3a1jTFNpSLFrgBPJsWwPMEwF
8fQZoOCZ7B2AdGcZ7DOmOU5ryukvvtc1ivY0zWelrM5K+6E37vaZSu69cEfNZUBcrBKVinby55kF
7JE9B0f7qf/LSvwAMkL9HCuyGaq5DWa5H9tREPqGecbfPP50S25lo66ZStCJr+ez1f6btlrS7WXs
c6QMToRBtIHX72mOUZ/Gxai5RvBZSSa1/9fFRGNBDburA1ZnpqFdVFym3En2IvvjpQZdp26dG/Jv
7/uqovrbXc/9PdIKki6gPLK31HMKLg35X8x/6Zl99LHaJjwIn/OZznb0G/ZLjSFnh2tSDU3yGXvv
Ic0MAa+C/D0Wco8Hhr5914N9daRBhhuCMztmoDngWUkn5rZsxzPX5KMj7VgehA4a2kJPzY2XJp2y
GH6ZxJMO5DnkVFyxdCIMulteOvd6IKyVOqN2VxBLd8EyBI5ob0tSTsxSoP1TpZWiF1wjdwtrJlD3
/UFPRsPeSHUkq996vi3Emen+VYvkig55jprNvUBPE3iqVr1eeegcf4mIh5PamXjzscPo5MHTWvh8
bG2EcjgzCra7kyX9CosMS5uiK9640p860+Ip24+Ax8SJEXeeFwThxDTs4QAIA9gy14+TG81iupW5
BBx5ZSgc4bsUv8Z8rbUTFqsKvPKxzbOVfbfCR7nwVyE0kpj/iY6FgHvf95KryrAqChjiJ5jBZlvi
tVGmA3dyqiqq2QLI5+RBzEGBETrfVkVlNC6R/bCIRDfHBdfAFhlcpYu+tEU5nmhYGE6HbPYovzD2
ipt4zmC7GESpquYbEuCAgc0mtYXdCid2UbvBfTU9PkEmTfAwSjjlqvHSkjqVgpgkFSEtMYNyjR1E
FpCEMxlL2AcEzn4EqVV1afUCZmFdJJKFOOHrDfIg4biMXprsKLSC+TrwJ5Y0g7z9iGoWAiW8uCjE
CMev8c86qVuldyqvAP+u2tPJlfjVHp0A1EA8xrVxJkMBLfqLv3sXPiwuZPvyByONjsAqfRd5Jil8
vrhmxYj0VRqi4LsScji1H2uYQAA5DxKvhrbRpbyZ3F7slSeyfMkQgPh66DL6EldfYn/5fjhQp398
ddZ7xcn1FnbRDFTbLVkOiEa5B40FGAtk4ZOkC6tlbqK3giXH5shk//mbDjzNgvbsnlywGFBBZLxj
1pvzMOwNlgQkGAI7Qogm7E2O8Q7Imk0lyR91zYMUZflAm+5+XHq3rYHV7M1mvg8JMQTMRx4dGP6+
Q0zSUswECh5mzVfgP1IvotQF0wbLWuinIfEmZT6sIP558j6IwfLkTHWeqw/hHzN+hBe3WGr1n+5l
YUui4icKG0A5ESMPHWvBm7ZwTEiQJ4jbyHUINSWnMN+i1aKr5vphBE3ndHO9yrSb7p6f6B1s/Rf7
f5YWgZwiTmHYdb1MxhVq0oRq9gNtQXOuCztd0zTHNlzLjQCKUV85gW0HnxRldSAIsRCYlFTwf3r6
wXjvjYnM0QV+XDNB910t/sI6MeVrvMriocuzsLRFfYbsUy9ZfEy5ZfOE0SNRiA0KFytup/VAxvvE
1LEEPFMCoc/ypUSawzFBWPD0750Q5OvustYtqk+tkJFRUnVjdA1I1wjs9/A52NHOufeYyDKHEICs
/ExX30rwN04IrwPliToYAt7uTHKFiz+49UdyRKloa4rA/L/BxPAchEjUMLwyItHISs5m3KbUOyeA
++XOeESSzdk84F4uBRhQFJDX5HdELVuZ8QmOGPX80OyIGeh0gVVrrpsvRqpCtexUZTkdbqzUvOoD
HxIYPWPb8dMDf2HlbZui7TUZC9RFlxz8iY6FaSs/K1eRRKUzclHBJA8Gq6pMhxnw0YSypOGLDxUF
VjbrfoSh3kJP+XEUXnKmbVLqVifwfjIQ0WMtWe77O5h9jr6MHI2niFpBkVIxsI/EciHsCPtqHcsx
K2KDM3+ah1FvNwWtncNOqO3TgAQDS5wkukmmpLMStqz6h3JDHdiPmnLmtOERg37RHECeJ4UjEHBy
tHVZCTQOtZxAwCYD+LmAFFw1ThVc/dzeBEz/ONoMaJTSoryw0J6xZ+TSPglAQFvVCGPP2p7zEaKd
O49Bd7gCbRrUXwT7yYaWReZpSPyorrFzMAd1mU94ArZq1t/djXjZ1BpZWdnRSlc8+3ERPwQwxwjF
h3LFET8MWkY94Z6NhzNo49XDijd4OXthiMx3gpV1wYwCCedU96xyDlW0tYZ+i74aKfFZ8DTfltYD
8BmnNovJwCqq4HboBHF8Rlnx/fxWd7/Yql2g003w8jKEbpTYhqOWCT10ea21OVA/56x+DklvdExo
YB3eQV9RFpZ5vLidwadEYGDWu8/bwIAWspBkOaixiyuzsDxd70TUt1AEszmAR8d32fyIiV5buGSu
SzyJ11jBvBkpLxdwB2Et8WaKC9/5DFB5cMXzGNW6vphnGt6NsG6hf5uEg9z2TT+ZcDZYQwtGyWwT
Ips4L4/qLICSAi/Vc5ONyW/6eCBsdUM/toabwPmWiSIrwSvIrXO0s+RPnMjGs7D9eYAsGPWcr3eG
q4z/mywlQS6x7pJUY00TJdQjQoXG8NesOe9Y06I7uSQhC3yi/RSu1LVO3JhYzHdrppyD28q5BoFF
nJKkAA/JFnDi8IzoM+PPd7IG2hRDgsLnDRYCSdQBd34Pd3QWK9rqzz568wPBts5zFAGcDmvRrHo8
XJI4VukyTOVyz0uJzQvOx9LHo+6DFkEl8wwXOwYll2UMKl6VZcJirKI33sbqXWLrk/hw5pddr+RY
dLtj79B/AUD3aJ+ZrbufVYgDB218Ty0mYmfVOzHJQGTBXr9Qs3RD+K/GLFpuPK1Z0fu8VeAYHBlI
w5JkaYcWHv4qkRBvnuZzpxHnW4y6BDsv1w3c4LleH3UvAtTekizWqTtzn2BC61oE6FpGEZHy2ieO
b9mzJ/tj1wCupwn117h9s0khPlNym3s3zLP1h+ZGXB4SUL66Xz7mURD57zw272Kw608nAXSA0MNC
IrmCizMayohDH9jiVwXp12cQh0aX5SpCmOOYSpannbE584WBqt5G/T66BiecS2Z82uYQ0U/AJg5o
V+pibyeRd9em1Z79dX6jDwvK5mFMmaIL4heY6XPv0AzqxTcpVk0p4Kq+3SJTNi1RSJ9er0HnUqZu
2lv7rOpiES1r5/PRsdV0rrSZ9nCCoHHZqm0poKGUvZiz1uTykiNDyP9usvg7wvvwJk/VsVok0xob
jmjLFA4QqKL6yeClLf50Q8rDwo48fV5msGHfvqjDygVfdvp0h2oJp8Wrem0HVa3xEHttpliGhr/a
1eksA3Z5t96ZyY74qDji4Xls0iNL/Uy7vuy0OoNfHKU+ESUHXH8QnMiKHHmNEpciy3hpwelNEUtL
Mx7yCl/gNBXuz6IMcZeRcMWew0fszh5E6Oypv6KWCQd6NdaAlegaAhVLwviE+uLJuRt49NZZ+wZD
vqxpZjVJOxPplpizXYE6+2ZzW7RklUh6PvjwBmWUPl+eSJJ9efSGtgbBNWvwCG8BsYHBIO0BLNJh
UdFH65+Rk1d15IMkw2uP6bqiD+Sh6BYyPJnc7m9YhCIMYTJHIwB2F1LiUHuHj2vt9t9X16ZTAsf4
l/RE2a+/ahfCf6kcl4niO1z36HUuoQn0UALHN9ViWSGOLqLFAgutSgOXcfBSg+O3O7JMWCiWVv8D
gJCHLSWsIcFViGwSy09PXjmx9larYK8WJUPBu+A1aK2IttzhnT+C5fYmFJ05jlMLejiBGMrvKBa8
yx3pxuLHwrkuD0egdnbC7gp8eBhKkxBpk2mnNf0NybV+goLGCQ3oW2nNBRik7E8uy77aXoHGIwtu
TmEKjvOixByxI11IkEmcvk5NYkctQralLNm98uoBgXZf9SYhP57rJ6MXSg/VyRVLJDJs3V8hozZC
X6qx+Hy4pWPcOczT58Wz8kmCzK21rYdyOxaRtlMfsD5EWM65Y2dNkD2vL2kiJll8weyqmIozRshV
3Joa0Km6Tbjd5vgqrCil404K1nVhqV3RRhY556uhrzHGIddc3+D2wWJsxa+Ry6Yg79pHeG89rqJ9
W/D9XKFQ9rF9Hk2ckwUmbUrhvWcD5XG8IraA2VHMRAUd0RpT/PTjPJdymq8R5q/AbhVRCqzRu2Qv
xK3FqEaafwb8yjxvCcZJiFr+4ysippOzrwDeShfPhSBx0lLAYRiRd2Kgapj69UWp4i1enMGxdlG8
zVHgHoWehyHu3ohm7Ur/WLpPMmmYldXlk//uvVwrl0w056WlHohF3PpypBpZpyBAkvoXyKVXywal
VPlRqgliowiOoa9YUfTD/51r+mB+nuib6VyyVaLNm2AtoeIGaSR2Y8zBKwXnCnmTBMMA6SoTv9Ws
aTKfvE3GqMov6nZU3xF5l5Wwq0kejpr6aSAhE38NXwZMlyF4XqJRKTD2jx5yMVfNJrDXuXaHON4x
h2nIMxApQErz21mmWhsxVEUx/ti2fJITLLy76m5wL1DiGWYUZVH4312dKMIQD1HRW/Vqeke3dPj3
SVD1pZ6yr6tTIbJ2ZXgDMn7ppKmr+IBSu6fH+P8oIvwobtj+2+fvNpazl8Z0T2Q39XmPT6ylhuUe
UucJX9sJpXV7zNZKTs6JsqLn94+AjYUkEzcSbb8/cEeHb8sGISf+FmNYvSxveeee1cQupbb6LqeQ
TdSM9afuokBJ1VzUMWw3kBUHpiIec8wwidfo1IjgiIhPsT/jbbKfQWJzW8U2V4RGQT7slEcGJouA
GNSs2/VPWTrmo3xsdzxIxwizdGCREnIPetKjvVDKoB7AFsvtQ9QEbik5rOVgpuH3fLyxhEzEA3Xh
mWDTbLOylTCjvCqdkInmE6hGOKShJ3HxPDbo+csr1f9kGA2TRzIsf4Z96+jUMh1M54+P+HjWrjgl
BTGEXwZXP4o1A269bJVMEFF5fW07KbSdxAX5Tw9TwHQBi6Da1SLoad9/802c59z+IhYtrxi4CSop
id5hDtU91r+ef4OmN2bW5FFITR2G7Lyo4+p7xN03pLAo60aBA2M064EPkpGQsv3pKz1Qz+nfWhgm
xjpXnTSnUKP02282Hk9boKPkClNWEg1mJFAw1Wh4me6wwKjtsxFk3JfUP4QIiGuPNjp1fjDoYFxo
ZUQHOly4osHNrn3FadyHKhTo56eqqRhYp7k/RD3e/vsnb7B/Eee1f1yWz0sZjvnvpXQ1C7n+LeR2
bTLIykCvv3pkee9b0DE351w1xBnCPTOTypF/be6Rj9bS28P2wTyQK1u3KfUhNR9dlNR095TlCwnS
5ZYpnxgYjVkZ3eNpjtQEl1Ek6FUvmijvFl3K2kscs37EvqM5JXperrnNICrJkDfMRB4SvU12K6ja
sJRr51/fkHHMFVjmguTnCTCibAIWQQIAPCL1Idcduf+5ewQ4BMYCTepBBurZ+cFwhDZ5sNUsknYO
tIff4/3LBjaXzqHun6/+2Gn9TRqM7riKzBFBEggZCmlkaCOgTAaVgTBJpmI8dlle5m2oh/iSfzQ4
x7Wm/ocIPSNKIi/miPCm1vYYpFo5evas8LY9obyyw4SYuRQomVUKub2+OMBnaH8xKJrL3A6WTOT1
/z95zVUoP2beXIqGoijzOrYBrqImkzov4YPD9kyne+REvCcXk4nYcAEAsLOPO+1+KGb+5bqTVRJA
p+IXeqzDjfbLgZ5N40dHti7RMbVTp4Vjn9GAmS6aUMY5aS+KQNc50VyEv42rGFNn6Zh5T0zA9VUK
b3IaqTxYCUvd9WGAeNHzzsCHkmlWK1W0kJCGs+mJGFe1VzKiYgnRNxlwDqCB4enGHxwXJJbTFCc4
rQjnt21g0+QgShnXVYW02gc5og0nz/g1l+FbrNuxWYo/NeF4gWeSl3D40lLIvUPdx9IMvqvU1BFn
a0OE2KxnVeDQ9nSFHUUL588zNf1CxI9X22rxVqLa208jY97jZ4XPpVCLxFN8hchEkSFo7trF8Vug
yRUjmWdPiSx1ZXa7
`protect end_protected
