// (C) 2001-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
mRGd+bwqZ/4zX/mpr7G/uQ3s1ePwwfX3a3oFA71tNsL6eI5Mfoes2tBi4koa/v+ZvqpG2mQgi4HD
yiknaW69n8HKIIYOUhY2IxSQUesVMl2vuFv+i/BP6sRoMKiBlbKQAGnL4DOBru2IiYRZv6BIgqYf
nJ1P+F7quMMpqUBlOfUNZfVi1AF5erxCCRegqmfDRuMiSZy+vnov+8G7POMq3GBCqG5RWyQyPtpf
5hmO/9dGH20b+qqYpQuTHMVmplsh/ECURC7LVzHAcKCX2OFrGrRA9jc+hMMVDAjMK65jDA5AvOzo
qawjfns+B4wZraWCd4g3O3O1i09M5n2hDkDyJg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10640)
jBr81nE+jozaEMLwmDP3RURMhpGd2v835PrwjGNl5FSGMhf/cz72zEMjbI1WoSUFUOIy26I46W4Z
CEHPQ14d2pMmpgbDD0Mkv+BhH3SM9sEMxunwl35JM2sq0YTDk97zB48gmjFRuX0W/yEWGnFjHnpK
57WCqtSTK7RPSl/qXKtGv2Sgt2rLkEWTOdkl8OvFTirAw+YrXzoOJUJU0zNHLUlDxY3/lo/aRpbN
DeguLdebNNZUqLF9D4Pwk2MbIgfte2KXZfNhAX+TLT37WP+NGMHWSmR3wpFGdTrsotdjyg3SCPTS
VsevqTkvLCf/AjFi0XwD2nvYXNckbk9w5z9JQ1luzP1o1uj14N+ck2ZglgkCNu8HN9dtWvlB6QXP
0C8MaiFdgem0m/qNxHySXbvt2HQjHniPlIZvsOQ36ct60rwzaMjsj/6oUl/Q7iAx+tRFvyojGhUF
DS+TKSN+zaXtw7Ttsm9QnCWgw7OWwcx/qdtkCGLl3XI5VdUWyFCPb2M6EQAqIKv0iTB8YW0vKxFK
m5ynH678xgeOycL41ETCx8RugFTnCnT3IA2D1zrlKbSxwb1HylRzDw78KttzftDXzKV6IH89b/RY
z9k2aISH/gCHp3mXx1B/USr37tdFkYORpEbjk4uFDrSp7zZXTpXFXwA0ebLCgFBpqJ93UGg4kcu9
jVPA3AD3Ns5GU7AYEMT7OWvh8QzINXQ8S9MogkpF7pmwky6dYNdfU+xlFfMBhaK6NXOaI9RbwgFo
lFRCpZwnkJYHRvPjNG8wSdYTHwDDUrmiB/kY8rVRruoyA15axwDPz5gSVqyMsDmpzG3DR/0PNWff
nhQwoKP2Ix62oyPwdqAyKa2k3lGwa4fCMOu2geNaMWyLONeVQezyPfK3zK16S+wdVH62egnry3bl
JkOXLgpfMiSWo3j5gHl4K9pkEI3J4gLSLIShmDr2AYh1A5l2FHZIgdEgjyhC/li/2cpD/Z5f4aCh
pldHfd7Trk40W6uSMBTXL1q7NDN9jfLl5wpXgEYPjB5+AHTdkZC8TY2WjwQKw5JypCZzjCXor1df
vjCpWWm76ahUpFp++FoXnjAVl9UYOXz5IR/C1mbQ8rEMkDF8GxYzn3lc5fVbQRYjQ2hs8ADQ+8vf
WxJka4NiBYHRDSFs7lNk7zqzsvIXSRjHkgYeFKwuRyf+Unzur7XgtYoy9NLixde4kl7NsibOFNDe
45Uja+NyNQHCqaYiI5FVnucvjRf+1j1bBxyNaNBq/SBAqLFYgWGnSKJUg0eS+UhhtjRjSSjqf3Ci
eflg1u3YcU3O4lPWmpJ4IxgnQSnMEzcjWnnzXDF/7e6Oe3XKPrkP88wVQj1Uu65KgqdIcCv/W9q4
rKpn8KOI8y0fMgp5VEQMnpxk5MC3dbCkFEqkeWGzH2xJLwgCIaOujx/JG2daA5qDgnJPZx+NRIjt
z1eqPW1zrCKEhZr+9KU1DsFfZBV228M54ep/HBQU96Uw7arBlKFKvYQYLOfUn8mZgZEkSEh12F5/
IbPDizIrhzh1y0PBZOumqji1lhF9DaYnAPkcwElQG6nhUMwrTbeW2mvh968DxCdMAseSReQhHWFX
fVP+oBqm6DY2h2/9rtnwwMM7uWHiUbrwaHtqLKXeEt7k3taKbvEyutJgRFtYqABALjXaiegT8oQ9
nX1qC7JL/BUxvWulLJvnEfUFu+070ogkRUekLgaZu/3NbxEiLW8Qg/3K3ccxGbFBb6nZwGP6laDP
I1OCe3WgBR2gqj76EtePFFJ8Jv2auiAA4tAi4Wslop1nXZKDJRvPELX31J5GEll0x6mU52bbOb0A
SJXs78C/gI8PCKkHODqSSeSXwuZIhwogsHI+0Sm8QTUuCncCtgXn5ZSh1uivl5JZdPji57z4aouR
Yxpl43RFZRNvRJIP+0mL52cyGDkUkg4r+Zr65QfYENsWAiKoLOGKmVRr1YcLWs5gSLYh3+ROUQpS
IlJCVx6O3yktPEqu8u+2HvjxJ7Sp/nL8pBpJ6liceOnx9J2x4WVnd4pGK+/xgEqyWLE+daZf/UvO
SPOi8cUCKlG14/F18PinqSlZUf38b4F4iH3pOUqWA4NZKyGcNMZdsXovVpDcZZniPP0WqXBg/vib
NgxY7KG/i+2w1vtIAB4QFJr5j5FJeu6GZ5xJcsZgyM1c8nDDZZPVTfgsFfbV93NLvEUUU/HWKHqb
9pmSISwZRTZrnMBPl/tqiZ6laFhM9dwtLHx4XV3FFw3iL/PVNtRgOFuxKZ42+bZDtGRIklM2I88j
0/R1o9inBuSpJJjKWOBt9PACVLQR371XQIMjSU3QSwN/idmm++0p8w73ujc1FJ65VuGfWIt4maB4
0F0SGhSKdjNnOdqFlwuYzXYqez/0U9ve25/A0AjYWMGvPvQ54kvlIbs8gjn/J6l3NPABSSoBedgm
zfPfn3TSkpUd2UTzyOWNN60yaQk0guhgtBNIW1KuQXxYWKKucdDv9Sqk4j+f3utRvNcbIQuiBdaB
GBMIYCnD2ZuNACwImpqw5ZzgdNUc3LlTKQ6RySY1ccnSWvxvvnVXS8ZtQ2JhZXCqI6+246s+b0n/
P7UKp5q61yXt4vDQuWquEcF9IksNTfyHU6R1YxfAlBq7QdlLe9grN8uZJE/ckkqT7buxZgh9yL3R
RTvB3+gPsLgiawLxsZ/aOKYEZ5eGf+a0zzATof+AXW9lu0kpd9snTKj0Ui0DIzuaX/BTwFd5+abo
YhuZgHsZOaHcqf7jEVRhjMNLcByOc8oiuBQOtS1Lc2DMqoZCPqF+oEF8tq7hFdVjrQ1h55fIUNOy
arf0EvaKxi5Rk6Gd7+SQ/B/JJnzQXEJlpi9tas0EP1IKHXJ+u48kHrhgNUq52WXnS6suo6QUgWOG
lYZX67cHNeSmflHoJ9DlxH+xTUeK9Tuyy02dbMffR1XYKtCWsT1K+No5bzBb56bm3lWTi15Pafu8
RuyZEeRoTNONh3MP8stxQQE4EcJHO+bkwt+Jxz/4Q+NZeM+b+RnQOMTKywszobhMmUiCjMGolXQc
cLQjM7M8VINfYb+rX3BkfVH5Zn63CJSyK429LY1HtwY+xhe/pA09nndlguH4TkizxL/jiY3qgLN5
SCD9GgIbe0J20vcCqsJ8oAz8+e09mVgQLvpRWinH/gkR/2vUqEKcuSYfVhI/gU3WS+7Y2kWNDWwR
6ElAKuzesLYCcq+0p0nqbhzZkcXx5ST2EizGCSkdmIAlEScXoTMNUFtELml8KoABRm/IKrJZR99D
eKrufbDOx5vqI+r4OqzMRwB3QcLyZzMieuIWyg6X8cfdec8jHmEBG4ARpRV/2DB2IiyzrDVjFj6e
82NjTEILBkg/o/pP6+gAwbzEAWRGC3IkazKYB+qyKbUDFO67KvYwcobZGdcEM1Lmq1t9NVL/G/4n
/nRyVQ0Y5czIbIw6N0Oi1CWea76lqGfFuRxLlk5jnWsq655ofyZQ47JfDIVJTAtgV6WsSX2Ieny9
4unDhJGel7ppS1ogPxj+LykUAAF09sC0+wnwqdgSxfGeiCzzVrD2OC3/wSOLTKL5Tg8Zj4iwqr1C
xVf6XNjQX9iQSViYCF92+kTzEYm22XpnmAnbhNqMq7iKO/HMv8BWZD99rQI53N3jjL++IoSTTrYK
BLs4C/jOriIQcEpQHI9KX4UPKCAskOiv6c2iaxAkk5HX8LdV5FvvF58ijCVsq+3p4MyzRamg2g7B
TlODa+TPNPLPoriy5lUOB6SplCKMJc0uuU+nVIaaKwAJwKsABNYtrGc4upE2JyId4iIfbWeeTaq5
zu2sW8epEhwtyRv94OLW1oix6Kf6tV3csWz5XPt5KgGtNNUDx18RXQwnge0t+uINSmNPq/V08/Y9
zDY8NSNCR1DoBWoRhWa4DEm63DncLLFn5M1Oi9aaIrKjfHFf3KRmqgkywJGqT/NjIum4GVCdTIf5
Xjm8rxcPSxk9GFYXU29OMAdxiCQx9XnUKLolrgJzHRbZyJdaSXM0QM+prC7dTwSv0CBT/Z4OQBxC
jzRIe9+2rUnTn+9jMG+D8Kyf5CoC3nOhgPvZXSro4S9R9C6bBQHQ2GeYbempgAX19pLGowxu+qAg
v2mfd6G4cK7t1Z+eNjOs0Et565c6jv8qb4qTHwBn5q9Y8ryYeiB3bmpD2afDg8oW5V5oKliEHwN2
GYstJk01o09R7aYSlAWSXgxzDcmuosHdsvzTaOFrtDr/xPXgk1TbFnspiCChXfWC/Kwef99hZGIp
2qi1Y5YrcrbT5n+YkEdlJOjqY1nTOUfwnrJvLI8z4EU2ryw/OSPH7kK8G/Ck9kKDaEaLuITYg4+2
V/0YAwgXCxJlJlMy3FGW2l7tHQU2aixyTS8BLrHSr/GjJe8OWnS0F6bjuzjU5PoCQmQevzOfpop9
M32l6h/AmUl+3JfAM+Askmx/bi+O29e8CpdlwHIEO2xL226EbTsyKncTCek0DAsPAi3Vb4QtFrQS
vi2OYTeAlo09v4T8uA76TNCu/5lSx6IGq+IHqoTvdUcc1Fb3WCjJiq0E2Fl5Rf3wzrOUgzKdU1fj
feknTvJEwQzUPXbn4qve4w13GDK5ll4+cX1tpfOM+UPZvVMDkA2i3n13MuUA2f+du4uAm39vts7x
djA4g6RCNXAa13JhrF84bPw79nCPklW7hMqRnNFUkFZXls/m4vKpQFgK1f8i5V/ofhiNjNokN3cn
a+GjiJ6bIEg2V/HlxOWFh6ir72iN8DXABCpQBM13IteiqYl58wAT60ZerC7LJC546jM1hHYC7VWB
/nMYH3FLOIxPOVToVYVWdwWb5e4j/FvAJ8U/9TIiY5H4W1fC0lipvuq/5OA3izIGy5H7e6+WdARE
OnHzOZ9tfRm4cuc5/gXsG2+QKmacjR0TU3ng1wwIUnYFD+2XuBkkHOA8ZmWcclEaWX7JXNnNMRhI
M12COArr0u0mjNxln1TZ2jzJk2IMEWSpMK/39ryUsU/LfF7wHaLAMjAaw5GjDhZhIV4mMRxT5irt
E9ZvffIBQnbxytEY5xIMofA/nmD0zXAmRTG++Zbkn/TL8do/mScGiZOucnIc6bVCVfNWZES1SEn8
wlS/FJqlizVwD2rhtEU/7hM4uZwF5MyPOYGAqDHjKxmMdLNPTCbWGlJGN2+9e+U1/D7j+WibUpys
3Sj98/lK96VdorBlbJyoOX0BjuvyQW09bGawubD/2FIDGo+R3LNScioBejkZGFMTpXvrSEKgqTyi
fmeVKI6H8dhaeOTjXZ+HcP3/NVbGPlJ86YsGWoLsprqHmo1hbMZC4ED+fBhgEvFZ5hntOQXtv2oX
fJw2NfJxaumLl3tPTS5D2ED7M70vfmxnsXwAdCtAC6FJg3opqnDSqdZRNvrxuE/q7wlDgxdC8I9t
PzjXn1HNLZeP5Y1TgZ05ARhHQLIXYy8jG8wichChwJHFSwZbGAJCL3K3dGqfK/ySogOd5mXtzF5d
P/0veIVO4QPF/XpUQGxGzubb31pFUTeRGCBG0AEQX/KGx3b/YGkHjoyS+c1apZMOGnpLZ4MmsReo
FP+61WAfeh/mzW4Em4+ioAGTsd553ZX6S5uAH4zHSqEV3yw3XsGnPw1tBXwBj3kPFH2jP55hoiu0
0YmeRS/dTIfFDAKNHpMFrGg6UOceXnPgg8jXufJM6imYopMqJU75mrktBpAM/BvdJbI95PJgVAW9
3PXEmiSQpXkla/HO90U448yfJMcy9sBCsQmnfm8DV1fZOHBkVy6OIdOrsoJ0kkzZTq40gJQA7/DR
C4Sq1L6ZxWQeSqQmKiw18AEL1/xYuJuco9mucWWdVN/fr5Mo9YWfs2xecKKQQIAiv5Bn+Jpq/gvd
YGilXgRYlulGX2aZ0PkcAFJmSF3sb7J/o36jEzNrmyZFjTKrDvq7ONYGKLqdl+HZX5gZJaSsiSz4
o/bF+c+zY5H2L4qJ8QdOO7l5WidouyqPCi0+3qSgZ1/EX4OPm9MATt72sWehd3k6wIDAcfPj4hWd
jxwqtoQdTEJN3myiiYDwCK4y9QsrzxT5q4r8iN3P+joxPiLr9ursJhMAKp9laoDYL23HR+fnZ5nq
Y7eWFdaXYgirmZX/Ns/rOLltWQ7+gkZTDwo4XdIRymPU3E1WlbqCT1DEHSShDtg2B3VkzqaqaE/f
XFxBuEZb+EzCB3AMmwIBjktzaRkkaKDkMUKg1zT0XGYIcLQ8CJRKz7vxhDT449OjgvwJQTxm/Kzh
gPbvQsNXEhfB3Gvhnd5MHs4eebZJjE/BJE76QyngEW7jQYDzGUVBV6rFcU6uEOBOQuJc2Srf+Jx5
W2eF9PeO0Bk47CFHOOLnuVUZXmSybfMFOGaxoR7hbHPggGO2XDJM5QJUyw1+/SR567U6C+n/Mg6P
Svv1V9VGYU0vpuwPKHcJ/AsprTreNfO9mpYgM54q0PAJo/QdxcTnK27kkykAseuWHKoc1ATP8+3q
3d/AylAZKgbyYxHJ5l3R9aOdCK4Tc6t87j3A5ZNRDPv3o4SxjvM4LMYLhp5WVz5batDmlk2coW3U
+Fe8hWw2vE5pZfneT7lEbZehmXBnIWveVGKb1frTE+zcifefgpspsSuAZJQUO0c2RAyE252nDcT8
OUDtiCnJSNRn9WSorXrskohwqd7s6VDlRwE3+Ujpud9c1kKFP4zmKLNQ+kaPWE25NF+FUhlq1B+7
nU1afTjfkv2tvZYlhrCgVnQixnO/VcuQWzoj80NoXLk0tFffXxh/WOR/vAtkswHCdCzSHSsQ5Q5/
wUYE88LX1MXwZXJYc0ucOtEOnbl4MmzL2L2LTeezaVv8WfvasChxrZhAvw8KBrkYedt3cYYxvpq8
GUXVNyrx4b3oXl6ODJKHuaf2UJKYdk7daoNyeI86coCWw6i9lqUA+LfsrgpqxCUqfcHJf97VTk/t
eBqLQcViLQEMgjUer00krufqODk5uCXTgK+Te6afAZPhh2OrrlMo/mEsw8ZqrKlNDZUQe6BGUbBC
766SylEse5qDZctcU5BwRvFDqbkPDbNURoieQAYklT5rxrgohKjbTDJ7yodVcTcvBZMABbstehq1
l/PKYsWATMbtdmoJ7OtNlE2AObJ3VWrtoCggirRMeX9t4cLk/xnED+QnRhmQdlZhlz1rgQiEzn64
iGytekDDk4it05lQDfoeK1ROtDJAUzds76fbuRdjEKSt9obDzUuSVHVPsSGENuf5HWecro9sYNO1
QA12W63uWpkQ4oNw8Du1lUhyOFbIc/mVDuhgddDpKKUIE9rqTxLUQqy61LjKWjQqYToTgaw4PGlS
05WV/fO9WVLXfueXte/iQF6cqLxGnhMZ+lAzbYomDd9k1YPrvLy3OOIjUvTk9SkP/GAAL8AvYOG2
qA9AjlSm4bXXCRIGqo7xpVHHif7K+GBfWyNfooocFVsPV76mKB9ZKlSz7jvXQwLfD9fQ/ZvtSzPk
B9hnUf5Hoe1kUFILBq3xSkAlOV1CA2okQlXCjckjnGq73qaSdrfNDO6piQVW4C+oTICrpntLE+5n
rh036w6R1rTHu3tR0NbDOqojcQQbL7MyYSgcpeYzoHXBCy/Xt0TKtSWlLIWUVN+L/A00LuKayYjr
gcjuxK6wKyuJXkOeG24vrYl94Eh6x//w/8ES9z+gSJCO7o0cOp4+ng1AhJK1U+UI9vJiF/M1Fjo9
9Kaj+AhKJsRm+PNQypKfucfKgdp41y58KmoxhJzbF2SG1hePoRQpcC7PolCsmntBWKSQcnWIsI4I
LGnh7tljv/LEi1rZWy+AOT2dbifECAlRZOtJhNaemZv6HlNyFV8X/y00+xczGJhOvMuPr7PZOHFn
EfzHIgDw8wF4PLy/IdlPIU8EqSGBXfFjRyCG6JPNA4iMSjiqBaMUXR8lQ8mXhp7QLDD0AbwN7MKu
4/b2CqN75O/vzEotHFUzF/x+/JYPtw6NaL0NUbwP3by+Agg1RWoOEvZ62hKh/y+KYriNrAqo/X7n
Scvo4Fs8PGw3gDAug7uxPSCAvn6CRDaLM3qH5QNL/KMujwQOn7YPU/0lS4qKcVOvcJo8RDebDy+O
uAs8Ih3MGoBv3Hn5M9fr0z59jxVP/NbRtGQrKk8gd6g8luvw/DVkHOxsspYqDUJTeHel0rznScXz
J80TOyAZPls+lr2qhC46p3cPtJylVo1vY5UvL98eMzjf5wTEq4oaVPFfQ2e5aF9T/Y5Q0VgfEQHq
2vKTlI2pT/xlkOgEScRDbWiATYOxQGpv0NpzL2aOl06Ii39JB9FWQ9qGPMAQmizTcbAqvlLla+Mj
ZzW2pVssH8S8l8Oq9LSj00U/wekWJtNOdTHr/WUvF4aLT5CqxpXXr5ZpSQWhzMD9yjKOnnMiqJr3
74p4z0fnlQnd2aAXnivpNkU3dq70h2ePw3PmbTa3Hse/kn0QXRTMk4PAsYypEUttEdg4Sc7YEaqi
d6WRUY/aHV3WXpZUrw4qsLWMOZiNHkkYvXK4nPWJYk/nKSu+5udr8vxN9uIaMeiXhlIHBHpKKw80
tFqb2VjjDpxP4D/fHyQxJ2yZ39uPEU0dvxQ5op5bznySWYaYPmYwjdImjaaXzwQYbpGMe4LkZ8w7
2B2moTXkbVfFYX8OK3gFIc4uAfFZPL1wuueUmFK+vcGJffL95XpwTbtkaAraWPlF4YuJhtPXrkl1
aTfxHMSNuh2giYO6+zA3DFiPXw+7HMB/Z19Ol+K264tE2gZJrL3GrwcxzASNbjNiPOOVLO0eDwa6
4KXHAs6OrtcAGPkoxz/AzkvyiBD515BXV9M+8fTFccmiWugXoGQI2I7fQFTqwqMRq2LTu5O1SNmj
e485qvgrwq+5Gn68zKQgD/MH8I3yQF4e39Vqqt1G3ARqbf7XhGtsd9d0lqKE5a1aYMeb9GzkYfZj
nFgV0BSyIQ6+pUZfkub8afG23qYea7DZ3y+dfmTc9hFSdaj2OrlxHI5u3BFkOEeD9hXoAofkWZZz
b2ZdVbx/k08ah/uHqhwwPzXvSmpveqk7MHOnROWBNCGr2/+a9UEasvcrVABn2ZCofcDwRvV9ApPL
oJGdhmSVCLA2jTdhDnY3/IRg/xbvK4MUA5n/McrEYSY9OXtAuRkUKtf/E2aaB5UPglsRaF4bz7lW
zg65m6uriRBjMT+x9m0pd/tIPcV9Rh0nIp/RCOn7LLVjmvwoL/2E2P/ls/ld2k+HM+O+qGy0xqDQ
U1ra4o01lJkFBsZjHnztN14rVoPWDILnJcV7+BX/7abWhqJ2HZS4vj77LAd8v8Sp7hixsMdGIsqW
ZdPR6/SEWW6U5/HnmkJpNZlBxMVwexvVxVp3p6TGRItFMOoLfFnusSPhzGepvm89r8/OhpyFdoGp
qnIlVb+r1YozdAmpSUkzAu2pqPj5sR+57sv07VRsV1x2MWkrismPH1YgFeB2G0ayeuecN69ua00+
OwyTI/wDVXiT/JVZS6kH0pO8wqMDczOLFS/EeSNijw7MuVlKYVNXkzxWTsSpV0oadd2Cm1NvA5Q+
QsoFKHvXQGTPzfEK/kY1K3mmSnvorJGlS79xgb9KcR9Iw26debmwhO+vnePv+CnfPcJkSvf/Kje0
6y9GyEW567qHOiD9o/TGcVxBni+BShPnvm90UjRUAvVECWQtDoCQkCmEE2ksOCqbl3By68ONumAH
yspy05YbQ8serhapdDwYNf2ZicxpL3+llKh0WWShtVkmYkvS4AK0Hq+mBPg4ANeV3Ykij2qLXJo5
EZRP08i4Bx74QhFcIVuCwv755oBTWaeQcyKE8eEWdEnO/GBuLEu+5qJMsVGn6z8+VViSWiL9Cw8r
jrd0FwyYxtUMSESa7kv1ESuhQD6UW+elCEgjH6hmdxpRtfcfC6xCMLK+ngwbmX16cD8SlyhPrLvU
0Ex/zhJKBvG/SVBiracuzK58PzApu6iENn2oV6dNUQGLC2p/2MufN9cholmE1TFzvPz80C+wIqDE
COgk6rvAitg32Vxogfm9z5KD6RFFU89y9Ub+DgHDmF3vx8Mu0latDTb8325stUTYqrYu5Ij4Bpaj
stoXZ+Q/d7M/e5cPzLtbxFEzTmn4lW6z1yXJm/3SXjSP7iMpA4iJvCY18OCNpN2yO504iBmlVA2U
DFhdAE2ljmH4LqNfrxIrG7a6DVqWISA0vWrGz6qPvl/4Fg19v10czPvIUktQeagB5bgbiD538p4q
AYH9oVgOXf+V4OIn8TcWIgXZEIQA0jI9BEfnUMA4IcEqrv+stLIB6pVjKy10LZMC/yBW/jBiJ4cA
/0Ca/aENy2jTKSO2XB3KO12AjSTIQ5czCaxAaMIyDc4IAKVfaadvM9sPBZKwoI9aPcCC0KsijQrg
eyyxw7hq+7e0MqIEAY0cSGy09Sij1ii7VjYM+OYTnm4d3uAuE3YQ9TtE3lWhCMi0aJ0J+762wMl6
0AsFfmdXnNH3e22WInbFjCBlUxvrewPylidYFYKAW4GoPI65jTCeEyZf8bpKP9nyIupkBt0uP53f
Jb8v1fFpp1Rjyy4jtSGeHW99/AgkP19ZnNbMbzql5E/sS3B7XL/0f4xCUK0Ymq7oa7ir3q2ysshQ
JeGsrgxZTX/PBQshpvavzxiBEu+zXtmbGYfmN5J+vzmKYYiEsEDrdxRRzgV1JDoFbkF4sfvdUCRg
a23vMh9u0seDu7Qi2pPiL8Y8uWUgz5RI2NC4neWt7WjhyJyTq4FsI59I51QmHBrgPdOlgKGPYxlG
WnjxB+OLz/sYpNhNaUJZ7J2rY/RfUq5bfRSCQjxrfycwAIM541tRQEbZb/HBRhQ/8prn2tvaVhbo
Kf25nvdpCX+nSlmfFAAWGwarsbSYRUXoaA5kCgRz85zku7ddMI2afJSDwGVPCT4wQP/ZbjgiKPTL
FhSHv7DooZhUTc0CwLKT/FPGytc37sZrQINJRlorcYrLHbAq4F8hEPMb2Ht0V7hDNKy+8SX8jB42
44dNDV0E0nH6sPoKroaxAP32FpLJ5745hWlNWIK+Ljg74tu+782nQoUj85X//uboE7NdIueTiTA5
UFMC/vt8m6zLxSUoDbU4thk1ym4BJ53EPT2lLP2/oU1iBKfFAXinMwiPtXH1eiH7VGQwIEx/KG2i
b4Ismdwu8q//IGWYPwsBOlY4BIEjNrETcpL95tsUWCJgO8vLfa9pu58Oh8TZd3EsPSk+1D3nTeld
JJesCCm9XVsWXlO14JAYex+jPYdcGb5BXz8sf/vGZmpAVX7VwYQrKeOPirE7sZ0Sjx2Hj1tWpj9p
H6PN8ML/BjRI4ccHwv/8xaBzk9HNciYHOGxOcKJqD2hzk815r40R2gtlfrk0Ggd0UZRsTC5DiZoC
FyMi1Ei8/2oDPdhfwF5ONsuhfr7rMLwmXZdiB/xNJqTvtw/ivLVgEnyNrICtsgOxJ3EoGtrrtxTi
me+FZMWrg5dZOpUesm0z6RdSxIAwfsjZr+x3fdjlQc6ws9upnHrWfkyxHcZiNcma1kiPFfy6POcq
OmcQvvaPvIjBJNfLJbzM6n/joXLts4fWfT6Bv9drtd2azk2Fwpv3kSH7q/Edm44SYGb2Kxp5YNwg
TbCJVEYRAVYhtxEbeeWsSSj3ypcLDJ74/1tXAnzZVlTn4+I5ey4K6uvmcoypQnVHsx2UABAQz3Gt
oUqgrmCb0pUFua2rjcpF1ZmZuwk9HI9ej27i2dEHILKFPNucWZkxfBonCXwuLaj7kZCLoD99I1fK
3MWIJXm2kxGojHZA3iHutMFBzc/5k7U/+D8loAmTglIjYdVKr94T/Y9WzzO+b4WnIMot3JkoDUND
SS/pccA/Hl5ExDaW/PrDIvcuSfpc48CqfamaUrlrwPqtJoe1TojeCGLrKHIWXTIc32sopx0yl0Iq
WuPt58fvBuV3KN7hVs0lMPUVGSsO7SnbS5JDK0fhSu9gdPaC6LzZwJzF+wkiVn9OJnbPiyb9wIpi
FRLqzmqy0nSBCpiIydaj9ISInDO2goNGDriOn27s8MMBiS7Vtf9Z6JpSsriSw+ttGZlqo49mfNkH
36JGMTJLX1vWw8JtORXVfFpiwQfRcaRDQVg2BmJ2ZNG2cZhjqgdpLwqnK4Nu/jjjUGcNFexMhKBM
cfAFZhJUyCBeM3h+k5bbEr7Qm3QNuDSFxL7m0DJkZ8kloM+wKffAX7CWoA9Wrs8msZq2jhAO/P4+
kBJq6CEFdPCR6fa2HIVsVykwFW4HFYabJdPUmit+fz8A8Ua9cEZIw0vJSWE5qmcrHYGcz4sW5JNX
v7MwqOz4p3bbB/904PgGh60CvStEyLXAHj2hSIwByanEgJ8cAJ0xIJlEDhK8xam5OV+JeLFd9h0c
uc3SFJcc/kAq5E1uaTjra91TotB5/lE7kEFlI0dWVHvNUeiuYI2/YJZBJg/au9dfmuclHBo5ok5G
AGKl/+9IxL9c5f9u1GqiNVtdcZzH++QslH0i2ZHTjZD1BlTktHpAbh3/s/xFSooW6lQ/gW0NkKnF
SWbDjgH9bcI9n6Wx/VEgPdgZ2RoIE2gqmY/MktN092kJYDqaQ8t+AXcJR/tWuAp5lkDTJ1J3HLTK
f1gtTgPvPujPpuJG8OA6LpZ/0nl0ZQqRPjPwLgRtb1Obi83xLY6NUNWypJMxdhlAtNLU8e9oK6A5
cCfNpXOVMIwcDtpJ80NXAEe3KvHIhub1p1lfCyPWpQDomijQbPZsQwU5X1rduZkCm3738DhdANpo
pi3SCortWQDZsuK59Qcanxe31bpr8B79scJrDAdqtpuWx7R4Jacyzi2y+x4Bn9ZFQJ8A7kWZcNmj
r4cFeGjumEuPYF9aqlubzmypvXUC1vsU0gzivRz7p3jhhdhl/CynmNcv2LNwscVsVZIG0epdcgZK
Q26QkQj4l+LQrVJMSOhvZNbCvGAP/oR3VuuHLWAEPHJk1UOI/g5n8Z7hz2h4PTa6oqsBqhGMd19e
JDa/2M/4ulLChizMSw0VB6ckrH9gtcJSmQcA9ZtQz4Cd5RiL84pX3NBTVHe0L9qLGnd4UzWLo9Qx
pvNdpxOhzsoCXr4+p5Ju5YrAx0FVUOx4hhtOMKie0BGVkUFDQUTZZI6Um95Ve+62wdMk1ycxJLFS
xAmdFullpyejreACmzf3Deu1RRattQpCwMrUEFqaowoedM25i3f/4zqA1HyMS2mz69bIVIf8YDg2
cjqajXqPCrBUGch0H7UlRWEMQLaGngd0PwZhWUAoElZDKnq83nwKySbC1koFHzP++U1z3Tu6w5xY
gw0baOQNo2tdA7MPp9tehK9gVIo1i6yBYSXt5mwRfIzPCCTTYpqt4Jx5uTh0M10fEbLPSwk1Mt+y
nXxrf+qNzmuUHbVmEMe9C4yM/JZ40XkqDu9PLTZhl2w/aMYothS1MIASa+sROA7W68PMZ/MEmruO
5YWX5PW5VJo597FqxlMecKnkjq/rgtNxxPzr3BuSWt8/E0H3DviCqevRKfGwOpy/aiMkhjHvnyvT
Ga1p2dsLMIAa9Jwno6i42QCev3ngfDDu7cvbVBGvVnYXxuqcXgaMRdN8jwP7qoPv+OAD5+K7V8Ji
8+NQeN/VCFnUvdnQ48LxuZUO1H98sb46lEbsy4CvWAJAKRvaiUcsPiaGM5Y3BRyEWgsjWXl7TjQu
GkHW3ydqOmBMlVq/i5YalEUMjulMIgp9zsNHnHAsjbyeC89etFpW/4/X0/mpCMpyHyRjEUYZVGeU
CvHyEH7HJgLspIBHcemOzLLLvW1eHGqFIWPtLRkrV/yvCqCZHEkWnHnB/F21IBaOek7zBGwR8tyS
NoB47uPjU82cU9HYF+92m07rOm/hezV62nwc1ZsuRlE8ShYiDLe7kdX8S5XFpCAkCyA4drzBp9l/
5lp9aq0CpriOhhfmFDp4OLXpdSQ7yBJftic3YBN/+ykfGT1S25Xn84yxkH6rbE0vG9764ROGRCkq
RptA8AmOD07kRPlzbPcjbkYbJlRMiqGe1Uex/eYlSqX62Avrbnqml3cZvQiHJd/QHas1Lz5KAG6F
F+n8Zdkq6aNg+avq4bigI12NAjvjp0/U2AlmvUAAfnLBOXojIqrYkW8dzGSWHuGm7tUZ152VzZlG
zuOOUZd+nj9RBCQShW64kdOskGfLZPdfkgQcVsNj4UQe12M8PmNMJkWfnXlP8Mok8bGewRGpgrKY
nbAk1lz3S2fNvV1de+TervdCaC7aNW6msJlLB7879f495kTpdpo=
`pragma protect end_protected
