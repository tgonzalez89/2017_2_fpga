-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Mo5pTY8W2niNd6YQJYrT4dIKljnB6QsjcBGtw8OTQa7VoBHq9EAAYrv5ygGUC1sI5a0zXmOUj16r
48TZ5DjVbGghhTNV3RUrNA9h0T/eWAVLERNLuf0YjXNxc5ogDnk/H/o0RtH8L6tbNmujvJbxaa87
6/q9oZ53Qo0uy8MlA9Q/8RRABnTRC3wr1z+XQD0EMioRsQHLQXRC62yk0tSCQmkVftjX0TZcrt/j
/9xL8IyTWBrLBbmSSD4XHM5lP64eB6uZxSQrRdc2YeJ095qHG2z0eTJcw98ncZ0n+TS7d+WXdtew
2zFWHwNV1u1v1SsTrBfsKwToeUUhxBrsUKrtNg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 33248)
`protect data_block
pMCZuaadh6yl7b0/TFeL75IjbcLHeDd00Ew+s8p88Y5o+Umnxle75fO+HkCN62kXJIDfqUDtGZ28
zBaE/ZuSIZYvej8kHgeoDJP7eOl14ARdN6aR0Z4+uv2KRWY17efNbXMBK/DNTq0MyEtXxwDWKHzN
O90L2V8Ls2bJF1xAWEMiXA/ouMnP6dm8soo8VBOiKrTu4iFLd+T9/iPLIDPPUmUTKoCph9KHWNmM
XC/3jbjzWKOdndeF9wrCAbIZvYYC9GC6AyMG4hJD3dJk2fQyAtMr4jru/c9z4tFqvXxWu95gZJxy
PbNlS9isXXm6mKBn50D1+JHUToz0DgkkI1eKxUaWDsWyB6FBGJklb78k0daXM73+4De0tP6OmfHk
1HZLxpk0Jfqd88wlRJxwr47blN+5lyU+5+/YE6MmSmBZCwF8oqr1az0oLzC7yg96R7icSgJ1oQeM
mtC2PxnIiRsaUPrwrnyZ9/ud8H2aq5uyB5GccHVzuz9j/Hw+u75B5cipDo64LnP6tbJ80hytY7PI
UKQ1neEXT9TVCcU6Z6vcTAOVHwCgbq5/lldrupb4xNBLhlXblVvhml0eOlsZremdt2QiHVvMm5we
8G7FU4TkC+gXayGUebYXCuLbdsrluc0MlMPWo2Z17rBVOue0k3BxAObGqHB4+sL0KX186rXe2u5T
JCV3DS+bNkcawN4YH36uZCvKFgvqQI1HM5/OyMzxyjVXp3pBfkrjqODqaMEk6DSpcF1oahO1/9mC
ASTpZedtTRIPH1hipFqVxORgKmqnIvjcIbBiDy/ZHP0QXxq3it57twaoWC7/iN1B30dz1oxYvKEv
YgOLZ06gx+C2XK6pCp8KEsn+lwp4GAPEMXOBO0gyMBic3AeoIYkvOgIkiCry5V1ew2PKtK+tu/wB
MULXtyT4xt4/4efPud+aAA2l2VB7xWhIqjotGtkZpUVBNtFoEQ5E+opEl6TMLQua7cO/GHYjsJhm
i03Mum68inyjvS7+LEXPe3YrcF2h/9RPF1QNa1IyT5djxOmvpkzQlI/yVtELccGN+8MXIx+5q1JG
AG/yjDlxl7aCnyTB/JG/jBtAkvjGz3FzqCz2SLJzakOiMROmkGYpKvwIJ6r8sPyHNjGnFHbD93Sm
a5jdE2qq4MXmzWMqay4QttgmqetqC68Hqf1YicKC0fpOFOQ5+kiD8Nq3ICiDl6Kzpu3SxcWrXJ5n
N/IVp5WvcOnoeQjFhYTefq+8oH1oBL6xLR6oTuLjyaUJGMlokldAGnsjXI+YNicTiFRciG+tmUx+
ZbKSGL720zKEFG1sOeQx+CaaYJix/nJapv6JEXvGJcNDa5WowPSCkTfK4u1PxcYKEqdn9Y0rTsKh
OVkGvURQoMNHB0H4zhI9aUXH3ts7XUFkkPjkHo2JM1o1dVwT8XTjMgdwMrHoQyzif/SRJKoR8iiz
r5fOhmvneCS5xe1QaRdmbA2QeZYyhdTR/uGGFdthW/ijHQhnbi7guPSDVo1k3xbh5rcd25NjIB4z
sB01sTPeQK40AQLCdrIW8rNTzcTcT81rCsLZS53AeIrsirkMlo99elMCzMkFxjwdFMPriI93EuWc
rtOB4PqNXlhUsSBA/hgmH/ZRTFsFdZwquF30cyUL9O09eWlVunSsX0LyVA0PVCVkbkr0yyynTN0H
M7zQB5Z0qDSLkowkTkxOGLalM1x+743P+OLjGcQQEiPnD6lRyb9RsrEOGMOXGVZdXatFQuXu1dWF
ZjL05BrGXR1xj0pPQly1ahwlgRP0V85FPIjxvfNVrBpDUM9T8N6uYvshTQKGUyMW+7piFKDgiyrl
G0SZYuVcM+Ta40lwehIAvqd21dshh5kYQ3Zo8tjBuPpsbEEldO/30fKlSq3peIZsXYABP52RB1oF
tMCDWxagCvVba+TM0pFVzDSxMc0yczUlY0Go2W/++9Gz05jZl1QL/u2xDw9njKio8BAXmHvchQg8
dbkVC5DUiTRYMeU68FVQi48sEo8BhNvXoo9ndae6CoLxncDBLR3w7KV5KC7Ff+yDKspx+ZS2adji
WhK1YOV5HlZnb7fSUjq2XgQmRZctOgML3RjvNoRNNxdmAke0dx1CH8OQ9wrddBSPK36aTfV7x/be
TdVkoE9lka9IucLbGJBKNBDCnEZ/Z+mMgoewaFA/pLx0POPSx0Wrns792iqKdDEa8FkfC/BcKd5r
D39FliFl0AegQkYhsCWrj3IBrP5Nlk/+mFdURZR6anNJF7ZtcJpLrmIM71T0yIIkClBEfheLNuDL
JmawdK4rgncsyojEXZK3CErUIL6O6w5xSUcpLEYpOgxbdGctVLFpNNLGZEkCI16d6hr8ZsZq9Z74
NhybsEsZ40QzTDf+BH73yd0D+ws7Sc3OZhuLoa4VQ4lTLHNHmm1aRLxZ8NSZOgWBt1G0v1/gIGtS
vo+Ur/lH50/kL8uhcnyqIlywUsy/xYClfhfqA82lW2zPQxQTdKIseOgTXbpcpIuwaOWOK6muHOQq
EqWQt9iY5M2tPajZNVY8zIS2SwKrsLDWtz6PeChHEwjwuDZfBAd7LbaIq45oh6z+/QUdvnQ0kr5J
t+tjaJfRUg8qsEsiNuUcN40yG1a4y+BW+OqcJPYU8ShJUWo1lI7Yevhdmg3NButjBZQPqDxmbNhR
ImFEOb9LeVFqnzQIiY68yPCXDDkKqrQceLt7U1IP+DYt5KbJfaShm15SAwZdvXbeOY9DIGD55BSG
vHIadllHsVpdPNTSwAlxJ6QuEGxLMRqka1KbOsEL7K12Xx/a+jmP7bOXM80su/6odM7gQ3XIq9ua
Bn8hXhjK+PUgwSrgzE56JBbSVFViEeroOZMLsmWCuy8iUS72P3igix5WB7f1byuxutL/no57LdLP
2PpR91AOsoE23vejquFlu08TKHEr7rqp34bIuej+HfN3wk/xUk2hdrRINDF+itoAz914t7q6h5/7
TEode7ZlokDFn4lpENsGas1T1TWJ/R6+tXGsjvKh0pCBPUGcFeL4bWzZyKRxVWve9qfr+G4DAxcS
DUghOBpVIqildP0ie08RC4aOij7jpq7QlkT3wrz4usj3ArZHvgMsIGmLJcom2sdH+CEUxMIeXc5e
qNqcfBmBj/3LdK8h9ehtFIibcHxTui1MoSLAKZ4xqsDeUva+/S/aD4QL5IbHkIpibK4rXbEKtKvZ
A+UnMMQVEBHTn8WTea627OiAg5fLaiAevQQG3+o+AcogmM++nIEOo4JDkKJWGS3lwjWHJWIc4pn3
GrLBSQe7+3Oyp+5eBxDqhtnjNQC99ApUSasRvH6MB8CopyPfBDzpxPXYo0oRrJ/o9aQLccx88DSr
Kmv2V5EAjQxtm93A6kzr7G3lSP6rdb3D3PTQpZ+jFfCDAxVdeA8xQu7S5zFJW6xSKHaJrBwyGtTh
YZbkJQmm2MeyVF+WB6NTgh7YCe3KHPxAw+GM0IhW8/j5FjvfMww5OhRnrj2ipm9FTt0/5Eipap5c
NioNKcqKnJfpoL3VUGxwDQWjiDvs5VY8RRV1WyKVcvR9p9TQnzS+YSSLQxr2qYcnn3+ivI1VZ259
8uPt3m0q7m1e4s6bhEEsW3lrskPOZxaOsBFanEXNHn+n/xoltmbUPAMhD4JFCr9yFDF5+3PZBTGQ
G5CtF14Te6f7ZqWAP0ifd9KhFUpFXUI2cvj0KAe0dJuqsZqigI3MSoY2fjVUK6eqLOwchPJ5XD/y
G9I6evDUNH4XTDaKS+h/XUU8OsW6tryuItt9WlZndgdXLP323R0e3pSdh9Awp3ZXcZOp/3suM6aS
exOUQZUxYIyIOtlUCnhRCC7DcpJeQI/iCCOgeTDjOV7bqhD3MjyYLt7D5XTxJpJpJSmSTPZF1Wek
wwgvxP2BWpPW/oiX+zu9FcuP/M/ETXSG0ITguS+AytsRMYvS9uQgo2HraVu7AatLjdMKqzTHZqXq
Iskn+tDIQSvmLGJqBvsgTWnQ1zriRUMBWAQSu58z8lHNoOX1KAk7bU2LTbsuIDbdNgBAhEzo6YwA
Zti5bFGxrMhKosfXXuLGr/GoQ/t6C9KRHb/wMZyCpxhjRJOAoIJ7juEXKWJsjS0SqBjmPBwWZS2t
WUUgPPWucif+g6m2fcisNaWOt3ewgG3ph/jzg0XBYGaWPP1FhtLw1vX1nX4Siz2+J9YrjT8HbpNf
uSWcEe0BeDr9C5nY7EVpPkIPOgSJSvlAyDaNBrh0qv+c1DsqLYuKiKya+82K6t4ADx+4vnG8ZT9C
KWs+wY4T51gmegcemT5VL0n7j1wgWXaXh8K9IWuxzAVBoFLMOcJNX5Z9kVVbL27oymx/bwPa53FO
PYr/+KJ0aqK+nutdzktxIbAd9cpX5+IqO6PP+dGMEadgLTIn+W+HYU91vUXXt9HfdcGppjVMPzVT
ZDg3JGhWrvJIYRY4jpjWGC8tqXAstK5k5K4exulxnVkHXNTQ/1RcaUyVpYlvQy7ThksQmyDieMzO
eqZS485SIQcQt8C5d6cDufScgv3ZRClYwsl9gWeduA9Lamh1ZEfKuR0bN+uBZdAe6iv0hbyDSISe
Esp27F9Xj1DsJGq5kJdV1ErsnbDB29jTWtEnLyMeIu8aToaQEwAavrnNgyGjEn/DUb7ykmZ1bB+a
5+y4DWofLp+z38B8abywRse/VqAi7xlaXYLaJ69kqIDOd8h8L5mEmTpcyFw+H/Z3sK0KMlQYLGqD
yQXTTN+dhAPhuS2RF3nlmQuK2jWBVc+4T29nn4Ux9l812dMusOy4gy4bwStx0XITR87qDeraKIf8
H8QtC98iLl2oBCvxkLOtBX79rWmDjIuCnIzrjISHPAYJdvXGOLrXoLosLeVy+sQMAt8QksFRkLc7
9jRP1LyUYiTfvbpmSzuhym0HuHnTwMvdi9mXkXA3Wqv5kvLRgMzVVVzyZVhOripEvJmPgapk7MRa
J5afM0FjphZBIEctz2aKmCHcxbtc/rRrhCTIuGW8fmq+jzKLW/3MIONx4mvS4GL50TP8IzTZWU+2
deJo9acIk5uLcuxbZk0pflM7tW1F7QAUOqc/Izlxy8fQTxkUwhb86Y/SBuoQITQIBmmZKeiZJ2CC
j1rTiO+vLjyCutOcQMPWtohJGs14eFPcULhvmB15DXrv4zpZDKGucI7a+5HBpZd1sbgeRRRVdt6G
Y/uvaGbX5HA9DpVcb2UTmOKUmrnZHzDCnKvTApITfhgkTtH117nhM/DB47Aq96qucBJQiVEBdSDW
ZZwRtx2i/aYgBdz0hURGjp9Wwt9Hp1sv4dJQva7OyIYP3vkT84w4D969pg0TPR813cJTmLK4mDma
YV4M+XlRvD7rWS5JD+y/A6JDLXTQve7DoPvlWtLQ2/ou8dKQ1jR+i1gmN5T0r8Ir9GYPLvFR51Nk
HCaGQ1X70EgQPc9Lbtt7KyF2zjRFymzYp+9iqJXA7+TZSwJYejvMgZ+OBw5NoDhA4vyXxJNsfUsR
n7w2B3niHFMR1mMIqXm2LDDYvFm1a+1WxQEOtboj7wZ3Vy2T0Od9wt/7PuZmc0vU8p5JLVMwD8Vs
PxTxXTyKj3IPGgjiFtNYymJTQTD2tE6AVqVr3v3/UAIkBbS3itXt1zLKylLcb185vUtFf/kLex+Y
7BduweXdlYKxOQ1yHKhJi8PfGXGMSw1z6G6bnBUK+ZGiYh2A4KNBGiSdB6ZHEG5UcESz/dqOH+rV
auTtelHxjkatxgoNuczZSw1awsDRB6h7vcyQjOroZiQk64We75OAjVALyhlhcOi/IFe6UpYbB+00
fadOM8hd8bjWZNvkmOULU44piTuE9xu+XIew0Pm7H2P66CGmbYdOatkqTjwZadsK1x6lEeZWikFF
TgCBY6JFIPQ5XIPujUzruZTkHfZimPeGNz2OC1oRBQqAOlFTBxo04aNfO1Gx0m2nsogh8tTNL5az
LTUDIii28opAF+UR8MydevTE54IDnJhdcmUoZU1cZ0TL9M/U3zdpTF45ZkZImmwi9apNEcOp9yKC
xDOA3qCfYHSuBo1EXszErBEyW61CIw+eTja2qssq4LngvghD53yWbLUbHBHz5jx0Tje4fVtqQtBX
Kpc5gJTA/VHUPnMhDpKplll05KwsGjeLPNS79Ve6vC/PqChw0fgIY+SM4AcL9ZW4nRaMzdrSUb+S
RDSTgWt6nOWW/Q4jHKr8Kd5T8VlBImYg+hKk49uG7BmAKZHG+0dBzbZfG5ItNxFN/emIZQjaxIZP
kRdhp4vZsr0KTfnNM1VPkRoK8Y/lyNyNd65i+Oon14xC6OGU/4itaWLLRje8Sga94/HCbGAjio/G
7d5kwLNXv92svl0M2YXGtQ+kvg/mzlfLG7Nel6v1pRaAWA+/6hFFvHgpfzRm5tiuMfKwXn0lMXGG
E/DOVxw8SaQQT0srLCGLs4iWfuEXLB71uJRHlpcfWHX46BWA+4VlDc1r4Y5B3mqCweKC0KEhkdgh
hgr9EDz9qa3ZZtuwg8552RLmy0RmN9t/I17ESGwSuq72iWEp91OruFPGsR2i6Y2RiMDLWj42FiIa
GWr1tr1KBGf6StcDmAhmlErNcjU9dhQ5ZElub1lQfLX8RuA1xZYUMfVzvVvIwbYLEzLMoy0/thgJ
Jy7rUL62ClFKoXc7krTW5FEb7nI9L/nbnkg5dR3jHVhsFM7Qe7BKMGKJHkiqC3NYcVleiN4Y33eM
czWXO3NPs/4NXke9lCWeNBAJ9tOvB8YxPh3PBGdDMLOXGw5QwBGgxpgjNxqwpfwIlaFD8fpmTxF5
FP3g4do+SCT7hLUJ+zUSo1lWLEAxV8G0mxG70tfSm2OLh6xZCWyLsQ86XRQuPBp9vFtxCBk6xjH/
60/SJgGdYaHiVL1A6JqHmbi0ephiwBzliaRdRbKCFD0S0fpm+XZCEzdsqAxH4E5rIET7GhcbWrJ7
xw8NvLGkYe4D9Jh1mxcocuLAN1xqNxsHKoA1xQy4hGlT1UXI1CuIQvYGuWWFqx6G8s2Z59YC+Elj
mNCFWJvs8F06jnL50xePWW36ajBuZek6PwFSJn6JlZxrv+Ni5zRkIwEDynJLmpc5f2GYnMKtYm+l
i4CzvY2pBxgcWrGuz97T67OPenwxGxUzTtsFss1LD5a1VVONz0GZY3/ptqvwXel9UzYnZdTAckn9
HbaFlxWNRC9sQDPo3UdcIStYC5J3q5I7+jvmw6M2vpwz5hoAO2LGIgBF2PHflcVcXYsGuPJNNyqD
cwCwd9llgLhlscgAMsEYX8OmfFUK2g1yY0VAGqG7CKsp87+i5doL5xPwFQbbO+l25s2R+ok0kNPh
2ZcNVJmj3RVD7UJuOHHp68LquDUQqpxDKsDnETAtTEqBaQvRQpI6qMjHpQw91047wPt+aVXvuPGn
cyyO0Gtbt/mNbt2kZ8g5EArhVAj2fbDGJYpCwuF9mJuxGRlju3fglDGS7m0/BC0jSxI94mxEVNu9
H2BD1obFvjoLc5KqtRVSerjWXUj+99FN8UK6XtbjycJXqOVVv+Gdm5OpjyqcNUpx7VMcAscqOVKP
+p1QKp+SiWckCjaYepllWcOMfZYhhLS1ZHj80Tos/SvvBF8g6YjixcdVbSE48Qg8AhpJfk6l5ZFk
f+2lXMdemhKTviWMoTje6U47n6LlGT4ysUaXumi7oZNCLpTgrjNaQuIvHof7cQeQhbu+rj6Umcyr
hIH7/PO6td5pv7O5bxfCOUdEuvjCZ1uOjTrAzHvdoLjtBpG3iZ68V5ZyXKcmH0KixvMNbA+YdhbW
VZYuMW3TreOnOYu+Ddj9ZLoluGJpVPPPUBF/mZ5zPptkKp9abf/WL2FWUVwhQGniCf3TEt9MhsAt
qYotq2NKBc1ZFSHW8cc/dd+njD/ytgG493YjQND5Dx+Z2neGEgvJyES1Me+3VCXZjjK1NV7dPBN+
QzaEfrj0iUydQyJSSCWLa3iu4dgeKJeVBwQfWIeIt5ac1Dcgz4esrNMaEK/ufs/cgqvf1JA4A/jZ
/lmVhhoQOU97Ijl5gUMcIHOo4XItZNnFUv39Vf371mSfR3a2tpyCEOujUNje+rS1cwhUUdlF44yd
JEGUh37F33INuxmmViJWgpRDNkcknFp1cU9Rf9aJh/33SyvzlXYADEx6MNF+vfZT/XHWx3sIZCBX
xnbs4lUhEewcBLXoUhsmHMcQgFF/ZY9dWSHoHnKPF6apVJWIGv6gzKBzk/WEx3upvU+KBbZqWOC/
kdqGREu6dCQadGYlhW/y5mDfG2FHZZaKHqJUlaXtQKc+7kL8YDM/hljc3FmYCm6Ym6Lx3c0alfgN
TzXvluhmaJNrfNaDhc5PG6zZqBbEYTFn7MbLf9SllrP5c9uuYz2HoQXGmNpcMQS3+nAOxCBUbE6X
9DZXpUYyKlN723r1HssbmLIc9H3uTDBPc+x+53vSPmo/LpIaFg2T4oleojP2DFh0eg7R9IEGgPPK
ecfHhussvXQha3AlRcGNdqODomorjxLb1JMLgEdnW8yHhQ4O7Cz9Us+M7KlBMeEGNeLbyizTkrOG
nJqVcSZHnGiCeg9534ErR0sROD7hrHcwtQ/+LZ6NvhkHLjRcZCOC99nDhS38G8Y8mNrZyPOBHtUU
QYsjtBoLQBYzyEMVZVcB6wsqLoEPw/lkJ2eGV2EZbJnH8TQBkDy0VvhxScXcwgvdeWWYMQPmOEUX
ZKq/kL0kxyegO1IMYP1KIYznMBmru2wB4fDtUJe8THW77ieEQJMGIFo+ObF8zWsSrzNCCvn1BmkB
y+DMFuBRlbdF06PUxyHsWzQbx/rLKFxuMHQBxBH7uIiuA19Ulz4rUelvkE5txcazlY573EeEvS/L
1eKAKrCT+NMn+WWyyYkMSNtIf8VHCesRrtET+S8QMrd0TJMXGNB15S0I9aVk0lpLRSYNYwnuVKUl
0UKzcO6bloAXDIZPtZqRVv76dbWGAT+p7WzndEZTQbs4nf3GAU6dGbQWnVtRZRfxIUQqgJBbd2QH
Nm8ijAogXZZP7mzYeSFjDPfg9plqthit1ccfIIk8bItZqciR3sTPZB7hmNbHaT8a8S+lQV53PgzW
ug9IxtVZ4jVwNUP8QYp2PSFg8PkCrTakORaBKV1XQBJf3pewgRYhtJnCoLdg3xIjDnLUi6UzAP/w
U99TS4120p6iJDwa9uDfZ17L/bDukQ/Sed2RH5cSlj175Dt/Kkx5AjWO36QCupEQ1FIms3j7yRwr
LHFMODNZc+Kp/anmbCKjw4d2CkNea62psTtFvvd4eDeZUyZDXMCEwD8nLfmvCYvv1GIOMBwk/GH+
V2K+Yk4PSelcHorPV561nz/+bw67qIuzDsr6XWDb2isKqgz7gLgBY/VMslZcLvsBemqbS7CuBJQC
kzWV1Eng6mZntcuGJY5EM8ktHsXAz+GYA93wQGXC79yoXtD2vADUt+4y9rWQdDDTSViW7DI+T6nS
/3SkluR3vehBJlC1XOeyZ08OHacq0lMwvcONDf8s7+1Tw2I/X/VW6f1GPZAG3g1RXG/NQaiIpTyj
E+ckH9QarPoHfJ9ROoXuIXSpPDcmiF4MyrBEGKK4XQn+3hpmpXBoLcb1ucIpR4Zbk+c+A9cOFMl9
G2RI10GRytxOk9kBC1IihWCBm/U0+zaVERIj55VxY/FaxinGjsYa72KRusuQZGpNTRIvJOUlpKqX
UZT2rX1kyijAetsqBkumWNz1b5LoOtSfWTEXOBtaGCYOWyGPTfIIrc7IP3XJJPckerl3V+uVbKyh
ZVNsl7d4p7xZASxtNkaDdW4Bi6zNANRZI+iFAf/9UrU1UmAil+iEoe304ykiza5uMLW4UPfwQfNz
gKr+3cB359btLw6vk7nvNv0MuHgqGsa8MCAQwwqo89zNDFdfJXrDzLLvestpfVusnVjgsy+awBb1
YRlpD4DrNSfU1S1e57t/ppsRpECa7XWBN3Kfl1PtiWFGkotNDpI/TSoVRkN96dmA4m5AUIHo6Y/2
Bz5RUy6t8/dV4w6116H54t3OsYvPv5ImnueNB3XkVG/y68XDXtUWZDSWVOUXTXDDES9xkxVUe3TW
pQcfnRfjZHHFt3cwuGUmtcWU0e40sYtX/dqLib+NuhLtEvEzAog3bg1Ph1o5GHMexocG7XeKLJF1
c2h8e6ELdTAUjcHURDqHpVHejka2IJfZ03H+eJwqBbiYEvtcQIHXIfuqBapmvRcjT4Zobm4gesMw
yoeUU0nFsqE09J2GCvBEVLYnY1L2ZuUrw6/wGgubMvAr9/+T5iwnZ1f6d/4nHGQJ8AuJi/Xx2rbC
rYYXPzMTDEUd5O6sUJYHKkTUVDNpl2V68JwkiAa4UNQeb5+xhztwhqD4RvFcuh8k7REreRvYf56Z
rRn0inr1YKZMhKbZFjVAbUqLZCM/UyAfOZN3aYOLs5gVCePeclYHiNZM16erckkG+RT3D2/l1QRe
FDL5CPEz7DaJxJbVWFw0v2zmFUmvh2SCZLR/NBSS7UI3i7KPBv/eABgD1KUZWQF6EVARh2chpV8M
O4WTJScbZyyIC/FKMRXYJyBc2xkolwtK9W/hd0nUPmLzFxzTAboM0CEzG1dPjCp7HN+WDX7xrSz+
b6kD7KlMq/bnuf2F8h/MM8JoFhPM61pewNlbnPDlkVH1HHNxbFLc+9LrS8Bb+VlfKaVId31xaE17
jOSZaiaNC4v+Gx+mgn2at7PH7HDlx4aBak6zqEZ5XuTSIhrGhdKdS7r+p9gIEb26/xBrDUjrGv2s
UHUni/BfWYx7ZaWm58ir9bshFPP3xDmD/qdYda2Qy/8vDo/LLAQfI5fhEbZFLyOKKK93g+4kg4ni
hfPL8kE9M67E0DnIBgkGWbslvSmOVCsCrNTWZ//LeyH7lQpazz7n6xiq1F/FUTTU51VzzhNrVjSp
sdJz6kFoUz/qamovzPh8TMm//jBzhUIOGaDTGPBj3jx31G0XsGs7tcEztokieKZhYdSFzRxjcvgq
uScqr8JQTywbNX1oltN4NXSxgctQq2RElGXJOWOjeBwbGDR/HqQtITtclpcU7bQG0Hu3zHcfq7q7
es7d97hEIMztfO19lHu3Dsgp44XwL3he4vh3Kla7v0xrK5C/ISh1JwHp+jEvNA4GluVhEXAiFMwD
22BGO+W9oCR8QWxqn0lmx9JR12JO0OaujVWZB/oFjn8MpvRyJLXRarOXelzW4yQTN/iQaCcRZoQo
PAGBWZZY/53Gvgr+WaOaA8Ft5U5/bXB75B8GecyVABcQ6ktFvKbA9GPGOfXrPZFwJ/cGsXqG+ntn
DikkY08/I0ak0NtMJdE8RtiTcAUdF9FjDT/CjkU2Sivjb1S5M47sgBZ6ZJ0LxUyic3lQ/BF4Duo+
0BxNKoSo/MA9x84ZQ1zfFmhBA5YToVS+O6XcJcOHAB9ORYkDhOuqYcMs7aOscmjchlUYoI07fxda
eBpnuoTaGndI5ajXZHtFHikUmepQhl26y2Ul/UGF8UPQJUgsrbpm+zu404WAAeQI7Axd6VIFWHkL
MTrNmXwmKfZFXrnsIuU/RY0fQdLba9vlnlgbzJc32+88NszmZQKNLX3urGi8bkbRPQw0oS7uNOni
XkYBXZ6598tsXf54oav15aNZ3Hu3wenFyhzkUlkaT3yGPbaEdskvkoh1vMdraEwP50FroigsgNAg
bBcWqTZYVBqiCIghWugkwtCQvOixe79t6+CXWYFwTCswQa3PNSRWajZoG2lWmiLNBgCzDWmnM/t2
6K/xVXZ6Jpz7/QFn53UB0mrhR7k6sW/aSP+3FRB95RzzWJSipDNK4bOWk/XTlBpwBI6D+Uw6ptPx
OuzLL4I/kWrcIxbfcH/cNbOXqOT52dZO6mOeFnRrT8MeP+ohb7Wapc3DBPQbcN53ZMSRz9Jp4Zpm
MMcKZjShsJ7SZGbBIBcpnYpihznqzdJy6Fw6CadQ38yP4RzdLuTif3eWJNXlJXZ9YlD6Ln2XqaMp
bR50kx1G1ibWUU8vqnt4rbrOuaP0Pp8heJlU/SCaIi0ovC5ZH+5axfBtG9GQ8Tg6Oe/8Yv24yyS9
WqfMh6Tud5MUJkhBcsByNRtgEoUA2bHlyfGbCjS4I0ClnDcl0VwqWqpQTR+DmTSooWM3EiLy5HRN
VFTY6Slexk03q0gdUGJTeqFPq+xn+gl0Cv2MlSFinUubmVTUc4gnDIYOjqtaV44wt1JZFNIx0ePn
EtO8nM8Z84SYGbPD9yYkuaZLTfkle1BonvoDrPBOR3Nd7s/dUgS9TX+VTfKdJYoWHVKi4TM3XO13
dutmUHDo0IqF50B+b/6Uu46+0YZZusguj6/dSAeqNDdFiYlogIpI0v1pfpn7m2ME6/kyPz8dBbZ/
F7kKb+snd0t+dJDoZmqegWbY1qnWTzdUTJGetyLlFn1YMBP/lRUUN9A6REM99vxA8Rwf4IKPl0PC
AG6wwzyJ7N9gkHpo4ohxEX6YpAXrKfo4wIe8cxNGdAyQ+AYDEOXMlLgXgu15RWulhcPod+Glyo+t
76nFHE751HCoPbDB3LrAQEIpb60IvJkTGQTteWvmzTvTiIJ9QCShgdv275aK0i9f6T1xKtQK5k4v
6Thf1NmJVvymi8wfn/6/CL/qqPZHEwHGRc1IlfJNUvvcfwVaBdP+G5C1v58rk9OvZ/KCQKR0Mx1N
CtPIvJNDtzNCtFneanwmg9RYM7OBYvxLfcHuk8Y9dgC1LPC8f9m+swSkuq3tWbWODg/yDSODYa3R
ShYhWG3UUcAuMW932tClDUwbTKaHpdtZ/3/6vF8RFgrkfkanZW0Y/DOBSE2XL6HFcJ5zWhDb3QJa
KKXxFraLQBgz22SCUORRF1nUlvVluVIMIht2WV3HC33j5BkvVC/ZTHydFTJe2PnRmFhPxMZp9zad
FUnysh5UIW65J6fPehlYayH1rOfW7q9+fwbXZS2X7nd/hvSkFCGqOycFU+JFBKB2ZootxWejrtYL
HTCLNLsMSO4IwLF9mXDTJgAVjKfoRmoMr/ib0y9OZ26N3B+Xaz2VOK91y/lqN5XubRT3LKAwquUn
JA5RCdlazuYovw3/4820Ya9wnxujx94193SMLPNgMUonrEWekaGA2ug/5ujK+AtNqrOLMnzIS8PW
DFnIqnuJBphkaP+pagd/8QTXMpdVXoxd5aq+CFmfmMWrGGH3cyokfv/M601OPfF8k2loTnXpTDNp
7/krsWn9+RWpgBgk3KhCoet+o68KJvn8bm7Bw6eUUIn3Kr7taLAi1I3wZPQ7SrHj9KGkw+t1z2Bg
TusFcTvXPFs2tjfa3OPOakC6tBuVFHH74c41/JJdM957EYGfespd3IKLRwWNLNTwfVXxCRfUF1px
3gGRbZJCf3fck0vPEjtG1Q1WKxAY9mb7CJEgl7aU8HPE60ryge6tjxmz84qOLpcuRinpZjqtKZs+
tJABAohntHYXlsuUvLu7ShDJfh8s9IQxtO1b24tLolSg/LdCN13iai41/LGSrcw3PhGuZzIHm2SK
LD9Voosr+CiatdqmN2sObJIaAFi5JWP8C9ioSgDCVje6+cccs5vGrxyA8yyUst0Nw1QWghPQpX+z
1RbN7IwlSrAlE36/W/hzdSEEnMC3S0/CTgkTRZRWku3GLeFfdcHBcX7B5PWzLCXch8WCizqNSHvq
6gwFbbrzpu9S0IuJ/wwy8tExi4IbRwm4kW6ecN3NE9Iz9xdZtVhbBpRVypimEE8y9o0RVc5Oa0te
72kGRYAJH3zwCCIR3vCdfe7ebjzBfS79QMOjEmVAe21nQQvNmy/LuqcOG0YtAACI1ZujAEgg2CpX
sAXzAQGw1x3LyMiZo6/JDCUBLd9xoRisBy01E87lFIkoF5Rd/k2GKM4uNCzuKG2HZKi2FLhUSCT1
gvA+KbBsqHf4Rm1w0L3GvuYHCh3hd199tE61KxxKQNb6EuJGg1vcWqM02TVqE2Uv9vH79Wzp+pLp
eiAI5gu/DgMPoDtX84CtRK2YmM0xEsDj7ymoCx//obgfd3hJDp28Ch90ceRNcfFUhZ6J+P3zYtG5
t/VkT1BGTSO54vHyFMnUA8OECpH+a90SEDm1CGmZ7vC74FVUlv4+9CYoED4aXNhRC6ZfMDu/yX/x
B1cAguD4XSpQFRtEvtz4Sfq6GhAduSmRWavoQBYWS2hCJ7wfhYLdrQblpc5xdSMees8pYZrp8xAE
zrt5xMGt440wjiUZeBSVEargBw0EeAfWsxYC3J7fGDPzAipPCYnPqMgOfyiiFCD0Bz3JJ3mFapVr
YJrepRqTx20wR7xZuBvBHAk0H+RbqdKP1ex9CXKyUrKXwb8ZY5dry550r44ziA0MqWe/ClA5+ul+
t7rhxJi1zTfzWKzV+vOB/wrY5c+P8QFohmVtgQC6r5Fh+wKGbiwrrCSh5lZmzZL6SoDWRB6cQuid
1IrP/H8t6rjqJvlOxHDOB52T9lhYVBRSUpensT+wjgCG/q22iPkn/L3BnWOBqfsB9GuVrCDDv8bI
fdiF4rq/gbdUlWUoWaN9ygYHDewTfLuMLfDEFZigaKHPLAvX+R+flCUcPGZMrI8I67s0HMaaW3bj
VS9JRd8TPynlJJQ5pD6psr8fSA7PTPcHpAWT7TPyAQgNwJ7dcdrBmwLgD6GFikFwgcameiIfeHwi
jZfDhSzX/JIbPCW3WMEIAG/Rh/1hv17NA4iz2S8igfHq6o+etSkyIsWvzWk2B5/iM+7FFCigEQws
aTMLSFUVHTrr293uh4XcL7/7W/oUG5XHhq4la41+6/wgo5DvJgrnfGEigbSXPrvjeoLErJJFRJGK
kJbG1rtG/o8ijT9vb5uJnVyasOMkYtu1ESzgkhHAAMER6cA1gyPcac7qRA11xokXobKv5kUIZllj
Kaby0PKWf+YZ3MOQbIxxeLvv2psQMg5z9FrexGnmat1jR+o0EXD0DxILrXYRtfgR4Y/jszt4Tdiv
1+Vgb1qO65yBpK3JifFwYVEVn/tCmVfO+ugyKCA+vzn7/5b7XQ7GL6FEVK1tUEhHtON6q9h7+xfo
AWADIYWt8+B+iv55nxcMW+LeCzzci9ZoaYT4xXsyVNl4yV9kIARWUPAbn4FsZz0yWhXqowCZtOVL
jLi78Z5qPpLYPl9jQVSohr0JL2jlt2n1uke213Xs3QvQX19LrYsMMVhOFqcD/LDiBCT2335B1sA3
AE29iR6gJrDnhLNTDYF1gtsB39clKj99EspEZu46xnBdP7Xo12XmwTMsWBtXIQOd4ww2iAJWtJFC
R5f3m7T7k+xwcV+xgXwzpUxK6jHtqp80GuA5aM/6qDAWiZmOgBUgmtrso/XoIhv6skz1GArwqDNj
wzyRhdzQOilMOz8pp2NheBRqzcRZn+hHyE9R693HuMXETnxsUujFo6CcWhJ6/VgN7mvC7sc5gdbD
tGfcLhzrILotZjg0Zvkxc2OmoMp1OsrRFLChzAg9aC2wDev3KSEsw1DYWVbTl9+IO1qZFNtzDo0d
mFZebPpdc2En+3+s2JBwOK878gfFtPpiqlNrSQyGMCs5Zr8kBKcMWdk4s+A4b3PZ7H/ceKT5r+EX
96g47BZGVG/ZZGrDNSDBvDca2rlBm8+pOhS8VcypFjx/cFJGjCfCZdk2MeQooT3A1/tC6NjnhKkV
9FHu3jt4OuJMZM01sQczzNG/BLNa0f7UWf6CU5j9Mdfa4OGK0SfwexJzAQOqQ7K5tHLp1M7o7bgE
fW5zfKjynWbRE8LI6qduGRu2UDg5d8byXzOrt0RT1gEanqJNL2nogXj32DPAaduwONZW+oCjajVs
dvSV9gyP4ooSU8MmMwhxQDcoO6UFgA1vmAZnEFDdgaEEhqFtbh6QJnT/Qcp5hojCV5Xv/60W+0wT
Sjnjuf84OxiSQ1+Ah3j3GJOaydX9h1C/0W6fGVCGO1btjXCZHe4FSGHukXu3FxbQL4X7SylEqFr8
O/9fv2vr+41nnv9nCNWTniRVf6mEfc6bbH0+QN63uNPHLpe29w6zfZvBhE+mKWXY9g1ddAHN9lzk
YxcBhenTp1R9C2M8dgWye5EDNVSydiQoLeEOK0xkB5XL5GnTQXek9ctjhoqu4qBwhaQkFMWnFhbi
o09hU3QATvSdIX+H2boffVDtMt+iuUwvFsAkNFkcPrNni3LNQMHndWvWOEBLQFl1jVd1H5ZtZpnW
5xQ6bS7QtgU5PsRdyKwbqogjhDoRRTnfvOXfoLgJ+boNHI32x9xV2/23KtxpS5sTNB/9pnbruWh0
sRU/3S+PmDEFfPoarupRU7QVfBadNLWuh/GVqvDAXb4pTxBl9qPIwSx+ZZr4kcpA1kI+sUVS1XPJ
g8kjC2cYVU/N3XXOSz/fwxm3E0EyrmSQkYveb/3RXnEg5lZkQM6OszKwI+O5adhZN+46bTwi2rQA
jbZJAQxjpnkaDeTcrOo1+Chqh2WNOSQSOnLW7YbCgcWaf3nz2+Hx2GKi30yIkn2CYYBlmILIeQbB
axCSb4OAETHovsV2jeqGT2ZJRTQvqVnCteumyskYl8jR2MywlA/+Cu+cGzmO4XV5wwTs9FiLfW1J
CBYoKn4irpE5CEJADba6wDixaoKmOcx/SvxPmsTlyUef1vIU7ZFoWKvBMgu6qXpW77cPue3+niFp
VUmoa29YBTcpB24EpdBXID3n5TtTxhaZyGG/7dFL7PhQ4xjf4IQJ5bMRZWSllz0IU5bQsfg91WJr
6n5VvxP5Ir1A6N+GFriWMnB82lIPJY0RoGn13IQCNpfLa9KA5awNwslP0Kh0DUI7iEIpCcYKKrZG
E37ZfDK5znSc1xS+mdYQE2QzzDS4v1V2/DV4aDt+KFlqHrUE+6A/c1uXwOydobRrKFe0b8MOOJZi
iFOG1oxy6MNbS+ZkWHqckYKU4sowZee9kLwcFFfsXDfH+s1H2boRspfqO2bfBa1sL+f1Vu2tO6Px
/IOh4dKVhB+IYo2Ng6pyork1gtGcOOiG67mNEUgE+/7vB11D2Y7sL3tK3AwS0TAhc/6u8v0NNUHt
vvaXgGkF1TmFI5dq9MBU56mHucLC9wEJpMxj17f0/z1slCSGhVzdCrDpANavh+2C75EwyKVmKL53
uDse1vTnvBZ5BHf8lMUAXKLF7LJHmi9yZMwRP7OgBWuxmWLFhQE0pHZ+poLfDw85ByYSkv4oQYdR
nB4EhCbskK1CX+Bx2UFU45MUDswYP0dRB/VimR3Jh8wfJbJfe+Ffxwic1q8Dv7Oea7wGCiYhW2+E
gy90rvkf1L0x/2LzYpG2+htO9YV9R4mVhjvUB4IJLAyQmKeUpMbNFM6QUX7XuGRv1FWWCifDKZDc
qPQRnQLb9YFbpKe8i7XXrIdfjq8T6D2i22n8/iX8FR0d+1m61icjgCmQ1zNQjIiVCYBshAehVLY8
kOWziyhWfNy4MIP7KOo75ywXcShGcmJS/1/fuGq8yyzmxq95OHRUM7ya4lojoYD7EmlgzK9GO6To
tz3Vx9E81q4Li/zhGy4tgL1pals4Rs3auOlFgtz73AVnDcUN0+R3cPWl1zkChh8nOFbOZBZTS3iN
O+ibKt5tIGliTuNfHDPwR8NcXdYUdMRXy+qApggpYllsUlLqBqX+6hHMrs1mMtW9pvzmaYPJ3E1H
Itz/T6w6u1ISkaCTWlXh3iaFP1dWVPS+w0pP0q1fn9mnT5BFcMiGM29R2/qm0p+z91g+8GFCuCWl
Uoh8WhCrQMvG4YlshJFosyEJ6I+bTqXipd9aZCqWoJ90F5vPRw6fvP1eP4wj8aWF59+zU2y56YdR
bCahh0JZy+v/PFbnppMC5mWFzjjHsiLnCY4MnKl3fMPDxhgW9xQtXdLav8jsL8sY0f4cfEeWHyG4
o/mJH5zAFY+rAcyHgjs89Ogvu1bB6a7wtWr/naMu7lUB/hpG70MUnIXpaWC6XDZLV/RGHd4Av8aC
Hs/UO6tKo+ociQP4jzRV80cu9u9bFvEsRfMwBGSl78w7wQt63I4GqiZHHWHHyy8XCDwTcV1ScETp
NmGoYgxUZzokvr74S1np7RSQCILnK6lq3HQGS2ml0mWn8DjBlVak1erFCLegsPMFmdxTdYcu0BUQ
zr4EVbXfrvjEMVsFVFARx6wpr4b2NtwsRr+jzFjg1Ol3yAiqX/6t+BLddqAd1Gp0nMge5js1NuF5
uKv8p9UGvl2Q2/deCYQRauYqxDC3zdyAQ44w7SskbDjjbPU5aedNxDIZDk589i7UtjHHF4TB0YMr
OfSXDh0nBn3Md6qKFP5l98vWungz4E0AfyEh2Zx/IBfkn5frbQq6PfVZcagiriS/tI54O+n0tSOJ
5xjGhu/YsuXwSi8O2Omq5YlJzVNd+N6Sgbx/hquqa86gCStFwGEc8P2W0LoBPrOp78u2K0RSbjuY
+bAWpZH1YCs7AADpB0Ugyqii1M5XkFpeshEcs4CkVmY2AiS3WWiTDWQJi3SmUNlemCUSCpWUm5yZ
zG3gO0Xf9ni6IwrQZ34pc4WRZN6GdPwN+2PnPNMAmBd7kYjyolazSpAB7GLlFt5BEIhfKzLLDVYY
5m2YportD2gmQF7sdB6npC+2tnd27OzkL2Pj0tUrYZ2gcmqoLd4kaN9CoCeRAQasg3w0fMueDhz7
4dMMg2UlKEKYvsk0+UgoXOKFyRa9fMZmtPPZFOJZjmJsVn7XbCaux+OqUwS552B8by7+CVcaMhbj
Pk1vXfb94PlnI/eyjJhULVWSwgU7aBwymW1tteNwKsipqXUMr8LlUO0gnjSFXhyVsOADncEjNhQ/
BY7RnCs1mN4jOQOzcefpxSRZL7jlfDU0BskS+oft5zQgL0EnCxbgziKKb8CQYSZF1GLLlOtp9utR
xBKTJ+sZ76Rf7KsV4hBH1oAX4CThRSHJ2chFkAmSqT0TxI3ZtgazNwZbdX+/3A2TvA5oTmiWe7l6
4a5puiCQgPJaMsNS3PhYUS3pV3ldHvwvAUoznBwsMG0MrAWscE0rCQQbwlWd+v6H2WuAru/DFxCE
XawI7R1D2DHrgztmJR4LWEE4bo98zvERcEyWJYR3pYqe2R47pKWstvSgsNf9CJhJgupgKOJsgHTp
Msw4TrGKwbjJmoaHRVYOURKBe6ptZ5kZL42Xweg3ixAt1fMk1bi5hLJW1CQewuSdLsQMN7T1LILJ
b1MXGlD2sotp0XrF2tMjgubicec9V6eUUwyrVSIXvOVlXVtqO5bLV0qa23wa+TO+f4ZBwL1yB0rs
O49aMnykahJVlG4L6Qvku8Gb+2u3f1KBvzyhYMczYC92nWqG7/ncyy5qIN6vxmr01JrBml6OUcHv
IRk7uhoDFtnYCsQohGaTHEkFM677djPfD22AcwxcAJJ0y0h4l/j1eEbf1qF6O3Yl8Tu1fKdvSet/
2WCowRCaJ14309P8pPIIzA5eRhQXEhPQgoT+YfytApsUcA7gSEqdvQP5ooEl/7xpjW4MZvD7zM0g
Vljma45I7D87oaNRwrgTFeIRWl9Xh9sVP6PJgwVUp+Ld2lLzFa1kqICdB2TMv+ttPlDdI1+qVfkB
lkGdWlxiunG3tp5TIbaBpgxYrpBx5lkpNTbByzo7zwraqxlT0U76Eq/x+jOt53FY5NvJiAK2SzeJ
h/RZQ+CA1XN8YGlDOMFZN7EhvmZbPW+/3nz0xOc4e1j6ZmYHbcgRNqs/OJw4dK+NxbzIcEqaQcOY
xJ/tj2Tn1SV1JRZqKvA50fJc99L0N5158ZUaG0LlOEABwybTXE4GK/L612tbLSURMVFFoSSE1oso
/xi5lZ9DVwyKBbWOBAFxceqlSTivuZGiuupfzZtkFjILoiWb3oNkEhLTxeKsIxUF5uvs4ImxyTY4
cBWtVhFhN2hIVRUxzVEazetS0DtypYqQjjJePP6JC/AhzpFlAPf90iWIVz9ovgotnkz3wSUfMzrq
mq1CHCnl2nTu097D10rWR77LHHVuACtKJ+P+HAiasIa6pNwQwOnZT4F3otrBYsYAcwcn+knH/sLg
WawG4is3SgiIrLW60L9enIbsiAD92+ogK/muM4z8vn5vN7xCfdy+yZTBdiyyLaEYHUZ0BlgzSAz5
9iKWWtE7DYCZYFEBcjKXfIlpy1iCcMTX9lS8QSBeZOZWNUNegYS4Mq1EC0tyACg730HoaQz1zj4V
YOdlqFX6JVr4DeYolvYP+Pj51M+JfvOD0aNjgQoXckl4sHdh/AU18fVD7t++uQq/nDiZVxAsj7XS
jUYQXeQTfeOVlRfeGQEn3C51M6AqOpjfM4t7uoTldMI/HDcWA+N3dkzOLxINGRfI76QfTD/iN1b0
GuyazLR/8w30NNtBpCWQAq3IK8akaJgt50NVDMeqiwi2Ny1HDzIgv3WQnw9K7DWoPL/jft5nAVRX
S6aWzo0f4Yc3RFgw9o7N/KThv9cwKWnBOA+l9XTulHhOVjGuy/JJvab8nnUrhshE2xiwE+Gw4EJs
3zKdmDUpeCmoLc5wVtHdZukwBJ4WsVhbwJdfSOkmk1EVqgaqiScSSYleBwv7xaQzlH2tEj2K3FjO
OUTjd4Xn6uGVjg35e0e8uq4QOM0WxH+oAjYMdRX0xiUyg4g9hmTD95XqIdWqlxswLLPW2ZRk+Uby
7sIRUfnbXMqAneuP0d+8TGV0iyYciMcs1yWVTSP0qKE5K8MXdJaf9M2Jd58+1B0Nb1YoBDEgMKsn
+56LPj3zaGWzMQyqBWHrhYG4E7vkm6wogfeIfH6NWQ0twy4FM/9R+nsrSj0ooyy7Mo2FqxN/RUtI
hOXF5ktPdifx6C5hZrG1cU4Ftme2narxObmgz1pnOx5rNoG4yTNJr1xHuxtyUMSdENed3V19NwCM
rgPT/5ZOFJIw6S2qVwlFYYPAC0/pEKLIjok0lQCkyGLz7f81XA7q76CtrwnKg0OYlBlIgajLdWni
q258iGsXJXs9Jh32YWfuaz/bL3fMvgWINTLYKAZSM6soEZ25bQ0rU7Y/Dkdy+IjCFO7NYNjbrNXl
uCFQxJQryzDg7SvB4PeKtFG8cDyOHbEZLL/nR27MmVFe4V5/dupVuQnO/gvMmJMRqYLKujT0h7kB
9Ndr6S+SLjxQI2c37OVK1IGPuzoEMoa7m2b0Go8YT1LIGoedF/75vwu6DH8rbx8nhKHzToSk9WOp
h1XiF/F7uYMxMNlSmz9I64riJZ8Yx5WKukG10f1TRvtB08shMyVZMaQYed7kh+uiE/zMhf8zjZ9v
RIGd853U2YCn8O90DCn8dRHqo++jOBlkcZYrd1aJ7rqmv6XQa6+alvWaeG2CJxKLpbV9eX6UBVq0
NFtkxv+kgwkJ2tbvPy+S5fI5itSNf1z542VWtSSnBAvuC97lDm3rkGTi6N0Ln3BCZgwmzwaLQbg7
w8bwjDYZuNW/qiDuXbbgWlwXw+7HMjgB7JdoccK+j1SdVOLWc4PD+t9EqaUgnE8+grPJ/qNQfyPH
u/WEq9ZDvS7qe24gSjxAt7gpC9wEH9XVSu6lNtRatwUbha7uySIdhuIz6cmge4PmCnFvZCNPS7vl
Z5o+iHBsQ22WxAS0wn+cUJXOphcGfuYQhxPxtNmyt1hXo+pBH/9eTt9g5c4AjJ6R1WM6gPLjRtRl
dO93RpeVtea5k7BhD4FwxG9/m279hBMu6aj37LHUa39bIj6XfKu3839mHBT+MclTdTIkVp4Gul3c
q0R5QOuIuvZqWxchGB0YFyJWzyfcmNyFP31r6hEz315AoitSmyYjDyZeU3Qtez1qkuZuIYmMz22s
497yYCaK3xjElDBFOMQwevlPvXKYsycP2oim9JFbrXJg1gmOuuBsTsktKFd3vitT8dAli2NB2oto
BtIlNB4LvCKED5dCAO9VKnxQ//JgQy5jDAaw0GO9PQQA+m7V2zayS/cbsphZAq/foPBNLjiaty4w
vTgEj711iUYPoibf4inGVuyD9BRDNonoyPwJG/UPwTXc4lscepEIMdj6Gx1i5BfBwcgySshzjNht
MBN4atiY1GqnG3nJpUOK3ODXfQ4VjEn/zh5ReW37YKu8kAunTnOvl63Omz8i8ejU1/CUpsHH8LTV
GK7c7KvzfKgw1ALVXFD7e6466/a0OPvk+nGiYV9KhT83/1TkJSMgkuylTAcaOko5Hs1h1SS076W1
cJquAIbKpgdl2qngPU42crI9fyGJnCIC457yS4TvFjtzcPnd9tRFCZfFvlqj7U7XaaraWEvQ9PdF
ykzfFTWKk+ONnaQxKrpU+ljmw1sj1QXgtU1Iy93BTgCSLwV1J73B/6xKcILmaIx5S0Li2RpCGPCi
9UqYHoxXrewwVAe3G5R5giPv8jho68BLGyF7FoLeFVD69jeooD85zoUmzOh3IohSY9RhOzqgotRu
c2R6Df72HZqgO1Mv734PTZCK+4TewN42hEsHGndVcbJHY3krRbKAGD0XTNpG7k0MXJO4mycr0GXX
bWkGQ2pfUR8msGiSErFDpO7JKVVl2mlm8L+HxzBqrBD2z4MkZ/DGVi5NGkN9z2BCifZUZQheF386
AZTf89RVjhQV06fHNBbGDtYNJYsYRr00+Icp2GKmh+8eulimlyR2iZzBt/01jlplaRe67YbZb6Na
tOczVrdCvpEWD2KFPQLeRZY3eR3V72hN37hMgd3kh5fNc1UcuU0Rhmy7xaOrtS2pAw1nwhhPtOsL
L45e+sPbnxiJEv5oQ4uAMEm/vUPABWb9D0VhoeEDbu06KGC7Zwel7tU5YuEn3gIt0k+5z4FCCSJB
el63BNRfHo4p/rDtzPWajpSWWg9fkilS8YjvOET5Il6qmtKLVgK1Ny4y3pDbIrqQH8T1wI7cb3OZ
7sjf+J1J6/RchaIcQ0o4hwgrthdLvAR0UNgdqUE8BVkEM+DG94CV5BWJxz0pJ6fW1Oa1PWmkgwaP
vrNQdO+IgXUb5RuhJnCE+rD2S0uu6EhS+h/IiqNpL4r0UdTXIDei5Q1nEROjkRF563jdVnVRUS9z
xADJeb0onnqC1BeL8RMIkYpSnD4UYEPDiR2/tLttO/nIU/5N8tqtcpsANFOXMazuwJG1Hmo8M4b0
rtDsZiKAKlQRqO5kFGZOcL7saYwAxpYLqHTlTZmbQ6Krcdtddhwg3cZ6OwL8jIq6TT8noV4W7ezt
/Dm0yo2dkrCnRyUziwK4ZU1WZMJpNzWZUCfJsGdb+p66KWiDBnT/3HjTYayPdXGNy97FK7OusW51
u1SZWA/XGgsip0DDcs5vYPi3YPU1QquYxdv8fDcHADc0GFyu6plNzAhH6IK/aRa9mx4RBZeMoBlu
0kfsOSUz+EO3RnI4/50tG80LrOiMK+uUN++mJZC4hwwlH/SMSmEyp7IBCFo1G3qPSuJd01HBeqCJ
rtGIplIYby2RYr5O81HOlynj7q99ZNCJ9GytDrmK+Z1wrNF+n7+hxmR87vLwRdypb0TAhU9KPCdx
GGfUvC7IWoaWuWZaRCnQwkRI8GAqRAkFIAAyvJWgUw/CsSQx9qlur/tIgKzUnHuUe/5KQ964sr/K
swwbkIoUqAaHoBB+906d8s/oPHj05LEcjdaGe7awADDmnG2DiONGWdl7Skx8j1t8Twq/JoSVO3QV
3VkvOoP7HPDkH+Jm3ZkA8kiyqVrXz5L5c6V8gsFwNKrlOzCFG3FWYzG2I4k9a28gmC72t9yJp0j3
6/T5vqI95+y8+cqaoUwgQjJaXvV5aLn2r2m9no1OcBuBRiyxVYBe9cp4klE5kP0BPGvrJYjqWaDo
RytqVJTo/LWBtUmS0NZ4Q/jd+S6iAH0ihU+CLlUw0D1Jd3OS+E9LuUGUkk9EvIgfOZiy7JmWgDoM
5CqjAxOfYGx47tnG9EFMlPyxF8AOF4vxgJuXwB7gRL92QVT0FGeGMXyMc+jeDeEV0drG64EYprqb
mx9hWwCXrMnnBuhadX5Sj7J0esUbZvLBqhntEPRy3qCZIFzrKSnLbhMjzCEEY5T9XztN4IGziyIi
M7AwUZ4icHWX06oxlfkgiaEzJiu6eNauLxTK5tKb+dc9BuOnAUUAp4l6WIiW8NI7T6HLCxcKBBWo
Lk2PJUJ37lgZTDoavZ+5A++YeyZ1fhlNAsJuQs1G82hEtSSfi+nUuqCZbGs/l/1F8jhNdOLeu+Kh
vJSblz+KyTpSh8PSkWhicYC9EClABwUcZW4cVSEiujE6blS3O7FN1ICpLKJ+u0jGT0clcNfqVWFw
SONjelz6IHsKsZFScIpLlDJiSGsMxmj6kf8Erq3T/dJLIeifAb7ZjLELoKNPBDSJuxRG1X6BB8AP
SL/H3fTaz5+dXnqqSi1f18zRkYrF0uEOMIg7UJBuOvFNy+oyPT9C1neEu38ABVvuktNJTKXskfuE
fZfOJ/RmetZCAMSh3A3GxpNZi7s50MQyTtDe6iID4DmiAXyejDVS06p84zat5eRxrCQ4Vd9o/Vcl
jDQFfjfaXB8QtIOOpqvjl43ESS61PEaOKynep5nBalHuggGbW9nVTS61v0hh0mmCanmwLGq6/yH5
Rutz6WMAdMBHZNDRineu4/mNbdWYj3qGYjfK9a+mNSHAgAAAvzvevHFrAQ26zrNrup16dNM5kiAJ
G3oTIdrththw0qkDPOxO5OSjUMj+3omP72OtUy+z/p44+CYOTMWRxec/FtzxKFvXzuD3UaNyQZr2
TwpFIwjBY+TK3uY7CsHTAqT4tMx6f020OndObewGOmhlKG15z0qaPUas5QlaOf0kRrXPtuaOmDTB
joDMJuuXVXul/Zkp7rdKv4Q4VZCEd5KciqGaC8uC4DzvMIc/K0X+pNfj8114+PtLwUf/PfaHNFgA
j5qbASInpER9vPmKp5hjRrRC5lDArCjiGdXIWmopbhJIN0Aa8yVugaRG5B4Z4n6eC2Dd3Yt5Uvnc
7JNNtQ3n9vQ5nNS5bAS2xRoi2uXy9lGtwOyAIiPIzaoqZxUhsKo7X9tOnWgYRul9MfXuiWnTefpW
Pu+RwGQfOr5R7rwaFhcDuHQR7bUWwDs1y+rwGIHvWGAjqusJR/n/f9arQzmAoyrL0BOfCB5waJic
u2QfElAMLWGEkRQq7R5OV7RKcK3FCpW/Hfbn9LxowD/tZ9RGoJn9rDSAzD60MGtXWdSqTCY7M8Il
3JVVXZJbUFWCWgrR55j1d9bYvWYr0QV/WeItE8mG/D0p3QCsLaZhZFoXN4NGKaespUiQX1sbXI7f
8/Veax1aPgNYzXCq3qHRY/51buD8FqkQUPAP+iWHJhoMknrafR+Aghn39xi17VtghO+KP5nmDZLJ
Pkb0/1QHHHqL9pxF7UMMbSeNAgBWfSA9WMW4U7rTraZ5gjjTGvTBWlpqMfMpPSN0iuhBtllrCBRp
Cjvmg2kBdcBhem/IK2i8q/9mtw9MoZKlvRwOiK6KtMNNn43VgjBfezJIiXWyQ7VKDbDTTPGWfgKi
WzRJFWQ5gAkmOLFTsRWmOYYIC2HPOh93WemTBbDru/K06lWsyl98y73hlwDR5RmeUD2kNp0KB3m6
GUdQ3nHqKEyZsOk5Q40iURuG3wYKZiQ9X8CrDS29JXlkwrj3/31v3hu2FcnndUGC3cgpd3mmvx1z
X0mD1XAPN6/oqiuxXgEEm28H/NfvF4yzd+zpz5QRJVFLboORtmwssULR2kA1htD2SnriGbKIqror
/JGoUvbQEEhJqnrrdAmLOfVWyory9bKxm7U+T7ObMcfsOZvpN5whOP2HDeiPS5BLzHdWTo64s95W
IcvHmX8Cye4OwXGJd8W1rVHYK2VYEPO+Rz//wyLviWL3pqfViXj7zj53en0prb1T+5uGU74UO+we
am+ZTWoJ3H92BlTSNMCXURk0yYppC5TkXhlNnb67ml7P2TNX4pv8t+npSRwajzWMdWr65q8aGFFZ
pAlHLbDH3UzTRsdKumSQGw+QruVPOYxedxHNWWzEGN8+dFjf/TEkho31CggPouxVJlvydmE+fqlu
e2Ooyoak4g9iR7TcFmzq9v8GcUUeWLhA1qYahJoXo1muLpbEvOwrfzJZADvXCr3YWcW/uTX2exw6
fifGglcbaZ9HN1B/J5CbKS1OjltUGVE7F40J/037DUidbIgat+zi//0LA73w//TTl5KCOyNFZSeM
+k0ut3+3dOdQgCTtcvJsajsIgrwBXqoVgrRNKWp0yDxL8A61bTKmwbvhypj3RoJf8Uj2VOqzlC21
gQvRJSukw8EOb/DsppfRRueNHFc/8t4zIMzYVHLudtB1dZqaFGBLnvRROaeYzIcuvNTh9JI8X+lN
SrEfn2qjTsAONeHvcZePuB4iBo9Fz69a5BAv9X79ZFHk85HtUitrI2UA/R+r+Rw9/EPrWu1Gmndz
3QdbSEVtmspVd3eBU7G4JuHl6b9vACoo3v86VygLRIYt/MGKHQyI/ZTnBBJphxzn0nVeezUe/FFx
YOTYs/hLKz5Nq8fXUSi83EHUnrc4ZU0MX0kQLKyllDSUAgO8QYDqfKGsL/asIhRaLpOfvAMR+1vV
T8lPI3YtzpUatfKe2sBFEHJZqMK1Fevn9cv4s0OiaIwLfq7Lh6GtkR046jMnbDzxobYgwdSE46Wy
2pEgF4597FiVkV6lhLMhv1Xuvx+8bVYaZmR+7EWYaKGU/4tlbhOYay8jyD4VqjKuWGFeHMRV5mBu
ImJ+stgH15TyLv4/ka9y7LS2Xse1dmP5luuzONebua2u4IJg2hUDZq3+Gpx31lRyJqB7+Z3k+3Or
Vz5cz5xIT+LOSPv8suSvxeR7IBY2Hnp1ZUxKJ0LR9Z7rG1EZN4V01ObAk8F5zutr7Jgc1juH1JVP
uOXQcqwxIwUqKHX/W+Y3FvFRXBlQEkI34zMLzT9Kzms/XaZKOn28JfzItEqgg6MMNyJs0Jl+gs7B
za8QVwtSN5cUGu7cN4xAQMbJiwzZUcG0iSn2cuXyKMzpaMe6iJEvs+DFZKMejZTMgIBaLnivxqrm
pBiQ/gHS7iDCFTWaVS0AgBk+RjElrYd8luXFmUOxyrNKyUwtIgkaMFF14Rij6B7pYCmnhd0dLJy6
XwbUDqwGBrDaW3niKScyVk1HcLQpj+cGObmLK0TITp6j92j7KXOAENYq4ToyMB8NO+NfmiSVNrCe
9CTREdQKDTKpU3Xh8f+V/LBcFU6VnfYiFYema0ERZQdj//KGFzsc8+9jvXuHB1naKbPk+O9E0o1X
sONwOZX+K/gG+5J8sjhR3seKmmhmMCIaSQpuNb7og2JY8KawT5ZI1+MRmm29uOVVycNDKy3uXauq
mLY2NLsXy8Ut5+G01Gi+oyMGOve/ZU57VNrF3B9qxQNl2o73LHnEjedGMSeMwuY3QehaiI5U2XWJ
rcxrAV52qT358FY/ABxxqi+kDmEmiuIBgBg3VsfDP76CzhzIEPs7p/tfKrfjDWOgHgTQXT6x7Jo0
Qe3GYKI6put3ltiqlRIQyZRHYwsKlNNnlaOZwlWpYrZTefPOrbCPrg5XXI3caijwlKi5MgYGCsTc
F4KFlAGAXUQi3gh42G0+T45xX+u4pqA4Pkv4/URURyzUJiv2L0fp5FUOP44bjRXHCVgSLaBo6SWq
i+KnNW0b6f0SOkCC7kyfMDEQ4Vpxnjpqp2vsTDfuJ9cIcJaiR6h6UludOCGSGsRCft74Uq3xPrV6
jZJ/bC2p6CVmkFHgPniIc6n9YY81jy/sEloahJtHpBcQTkjTn4CO+yELxhO7zfTefJmGMHfbazyX
1PqUr2nfkZX+kYo+lLvFEDZIW4EX1ITyTxQXmqLucivgGZv62sZ8SaD2M49gmjJl4NzVRzzklOJg
KVbbBLARrHx9taIRqZwGfpzHrzAatqMwm2ae6wpij1d3QqvVgA3PrdLU0rg9D+V5CHb39A6t8cvW
gRXLAguacDHzCoJP5QZBAASK9/GYKoIexzr8S0ilR37A7NN49VeeBx2eJdggz2oI+vP2/k7pAsAJ
Rb1X7rsWVRl3bfS7Yi9oA32YhLy/wnnkbpMT8jWhUee2rn8P5sRh4CxiYRCw1WyqScLEJKjaELNz
NB6QuxmrTg9ubi9mjuHAcuYmQiNhZMZaoH0wzKay29hPn3u2IEvnTsQ6poDo/g3jwOMcEERiBRNl
Izujp/r/FZPENLadBCRk42Jj4kD23bbmXrF6GV4VT2srmKeTj+VHoTtwuCCuTG/wH+rY92DPpymE
2+j2tJR89PBB/ma9AmS7ngDXBHz3zBa/wDg6nfzGko7zlhVgdJlUZB44rWWzrAB0IFc5pKfMgQCs
9lD9armUB+hI7AHMsiVN9kN7h7uJe1L5x1+v4KennqStLBLDm/FHm8bp+EUtf8od4XAzltmxQM7Q
KX9Jg/6LyPTuMpKIeJjdjezinawHuD5H7WQBwPf0NiqcQ79MQvRits2X/MywRaMZxmq1xsitOWkH
LX8bs5iwXBr+FBDskTxKyrC7uo5JtfJcFyuAC4Geg2sPP8S4AUwFnJExUVuZpv0YkDVt+6fKuVzP
/TixbjKWdazxh+cZXtgdg1G+IaKyZY2b6ueBERKxLDKWZ4ADnduUtdr3GFwmi5s4DF6FUSvKA7LQ
H99vrVF4E4uYgUPwR56vR2yoje/zQy3J2aIATiaLpz3WR6i9wKUuUPbLyQj5iSuTfoRbMh8H3rvq
rMjxUjrzjrb+ysOFuBKFV0KPvBMRQxt+KglFK17cGLX66nLMWAHz00oXK6U9YsGACaxcJwidOnLL
udDnWV+avbnHlkvWi6oyYd6XX6db5/dmVdjZbj5wHR8Ge0oDMh5q+fOw0t6icBlL00904iMGzrdP
N1skT2egtVqvGylDuiHgPXkE3dkzTTwLIXgJq7M2Olf2z0FytzMQfdY47PwoxU14FpluQLf+tvz4
nCyH7QEpYyxkQpZiz7y8tAXhJBhzG1ZfyqTEj6DxzVqYrO9MmxpuQ0P0Trdz14YMIgKH8T2s5hM8
IHCfT7B9daLw/TfSbxBqmQluMYAmD5oVbZ91doJSUTMqQ5daT0Hc7nSwXx4ToIomDA93QPheYvRi
a/a40eCvWBMIv8HlSNeeAAmZlutSxzDE/o1azau1m6fTFNjhdWWkUa1owSxoljXmgHWv+YZl2wUz
paBbDTFsxT1L2OdhCVqV++GZeYszhJxnZWHbVXzyhhN5Hk9wZoWjlaDmvX6WLoXpYeUoaoOWdg5h
kFW8XJqttfDI1zhTSSkhjpwsqpTAyJwZkjsmVUx4dx/N34G8E4S4A1HC8ycsfG15FjGaprPwtaQ7
lx/E79/5pgWW9dXMVQyyfjW9ytBGevVC9Q+rbgqKRvAjjcbjw5bxPXu2/yYr8ShidQTC5Qr9d+Sa
SoG0Rm2VkVPuEsyVb1xW8jjJLV0m4fjhcVFUrchb+YFwo5M/nnXWR+1ZtiB+7/plLxvJS+k+D0Je
yOoxey8v6ga0m+tE9qhwU+vW3n2M7rQ9bTGsXkdGxZeAT4dVyw8b9R+pSSk9fjW7R7XLPJD6lipk
3WVGpunYBHO0Qzc3qHPeBh2uXRSO/+cmRpd2V7WfKflr7VNgAdwq2kdQn19PZa1V2K4+Kr7ublvh
nr2Mu593MGMq0at4r4ObYy42naCNiNZw1QoEFLPSuRAr1kRV41Zgu8MRktGONYrzAtuwGYcYQvps
I0Q2GC7DBrT/CZoYr6qtcj8Nbz4jVLWJKRYL3ZmVCZYRZbTAXHsr0zbHNccGwz5+tu565DLSAPvv
n/euHP6egGUatknZ0GMhXAeYXXq7z4yf2zLlIriH3owkgnJ/p4Rsk9VANbGQHdEAPOrZDJxGSq3A
u/bXlmqvT3EHEQ0Mx6swHDjH+qFOP0RnzQVZKfilNvRAimU3iZ3rDsdxgI9mNmJ6WNKU0FPsBO0s
7BCpARBbwMdElvcL3wWX+o0hR3PoXo01OPpXT79Nyn02XE87F39bCzMr+hypzZJ1NG+ZmL+W3h5r
wRrNmZPkNRw6HcY4iqLGZW+90FTnjIqVcYpMcGv6OOUelQpWT/iumIhCMyZhjDHOlJXXxOBf5tqN
4ngc026mGm8uolXK6ktFc3KBYXCG5PB42HYdpihKsiSC0VxghmxPM4rDLF553HsgR5arhNSu+xs9
z+zl6b2ILRJoyiLRGEQVD2XfCo6JbRVPwFjgxKyHFpZR/mW0t1lyJYfhlFSa3L1tgBhTFcmWNaI9
8yxwd3IcTRTLZWJJXMQF1GG3YfJ9IN/oRwF1dmcBmyAh6bcpiZOpcu7KQAMtucE4hDOiZ4apFdGF
UCG09Y4FFuHVrQHVL5ROcogKrieOXrjV0h7mIbBsKaOp7+G05uDXskVW6ngjlUpbaWzsUyhshIIV
FbfYLhAnT/etGIzJpxVgRXDG7O/k9M1FkBmZo7afbREmdA79Yv4akaEGsPqo0WN+pCxqOggDWN0Y
vf7ftos7HW+oCDa8G4eFRektn9BUhVynGPEY7SxVrcluyc1CmBrWMHomgEBB7jPyqMF8btmzYMF6
UDlkn6Wwx3RKfKmZUT5qoEymAbtiXFkAlSooUU9YIXz9lpGeLcRG76IR0ka5Go5SinyC6lMYu5bx
Gu1KOpma3d0B5lV7+mMp/N30fPcApi0VuGWwuzsViprZrZ37CmvWwEgQOcl0h8iCpCzy/t6A3Xx/
afWNppsS09oK3yrtI2jZAg64TTdhDxYllzeNABH+8as2ARxoafjD59hPb//SAQv8/9kaW2bWhATj
Oqh2vTJNiZXYjRK6SNNBSxSY0LKJSrDC2XJfcP3sP3S1SXOfZ8kPbQnYmA6gS5Ugme02zvYbcH17
2FkpUJURxGhAgPu7oPgclgY/SuSk5XBo13Bish8wJbL1BNWUB+XiKIaWVRsXIvsGRwXBSNTmtIMw
b6Mg3EmVsxQJ5i/RM3mIWrm6MIF0y4ULeyTy11gm3QUz2Gj6vI2mkmqRkk3guq1QQ4lTUlPmRXUI
D16KrTOJHER5mV9ZTr0OCh9rU8pRNNo9QzVsUIhj59FIYU+mFFQSKvxpb7rr3GsdGVIhpMnCKO6F
r6angLTeWlk3wFPL02rsW1U/AAzfnmRAGadiftDuGPc8G1SyWO07Un+V3hZ0RXmbeibFmCfse6mF
B+Wnzwy0Kae4xZsr2ZiV0JQ/61GNd078YXEh/nDJdJzAbRU7giz6aWA+wWeZB+HTCAvxxMOUYjX3
+KJsGW6XKfn1vvIzSM/Q6tp0bT4ROPBr2Qq61K6W5GMKC98bGHmQHPW1yv5zp8K7Wb1vTd3+a5rV
qnh8whpPdttWn4w2JNFqb16gkZ/mkg1E1TQkeUARsKK4oFudy13O8KOTUVt1NxRpqNAYz8zJW9go
eGS0/Stbvqf9WnCZSuYFPP7DFHWOWfYDutTXTay24jWzGenHifaadjYwH/dBbGSgZPHdhAGlLWkl
lS9ltp2RBrRGLTFIpgpZbpMgac7vs+LKRB2Hw57BsoKReF8b+gydnHPitCCuePrESxviv57IE7k7
1ywTviU8DZBdsntnUyoStSNnMPODACZxK4nwmjUXU3V2zQJJhfT7Go7lIJauRE5CBgv4dkuk8m01
xYpGHVBh3w4HcciVCjCw7ShiyKTkSbU6e+oYTgzeC5j6UqPot1aTqTavLG4zhV8LAwzF0v6pRE67
IoF7cHVHOC+0tahnfQM2O4diA1fjuXTcIZaA6GGJgD2/H+iGpszC/zvFKkKG7B/Z5lA56HIkLC6J
WwTLGVz/Ku39tHrCz+Bxr/YdzEalUFk178tOyvGe8aRYFErzKwmMy+M6Hh75zcdOX53LXS6Lobe5
boj/h91RcGUq1xPxiCi7ecuMi/pIK8MyVddLj/zMB1tSiheN70z+pdqQuBQw8F7l2IGZLKnQ1S7+
RGve+7aQanjZpobSIF4GlVr2COD2VosxbgmOFQ4ge+J6PwocSnH2JeaHKQl+5vGvMNokMw+vjXKw
BKIUFdfe2Z4P5qGrHMM8XlO5SWwJCqrDxcnAEVWN29RIamXG1CdUEYARdN23v1OptEHggXHz8BtW
f8tU/5mVfBETdHnNw5YJnApwQdsUKFQbZdbQP+CKQ1b7S6nBSLq8tCy5v7M6NwNhQVcIzqSVcXoB
JQyz3yHscfrABdvhBRVrCMMP8keWjCuEZiPVJzel0FzSNTfXXy1fmaq2Gau5FP7L3n5x+R5YbNCe
8CDIc5d1+Mn5KDzI5d23AYI2AkMItT61EDqfAe60UR5CPeA6Vk7UwvKq1N9RzW6oGSEltVEcA2gN
4i1KGmjFPHnyrOpWXQtZLfl4h8/LBSkciszeUcYfWXOmYXvVEXNa3ui+xNFslQUPt32GwjIwVfaV
Bf8lKkT3S9Ing66/bGHEvuGTajjv8A9KgMLY5hVRT/p+ubsR8fxKrHKh7C828cRCBhBu4zBB0FTh
BsHAloSpYVTLhh1CgwPMhMgppKUzXrhFCJZR3iE8oRu7DnvpheWmlBSqeBx1DkCo9D9hh2HvPYyd
7TdIZzyEFX4EMkYvo+Z1ucWbLFjyasvYt55/HV9YYMynZbqNTwzfKqmaeY7cQRpySLXJSaNYX1Uy
ZyMNq6IOCnCT2U1T1mi7ZGWJonmPvz2lhUFTlAfE/hFsfVEmsSz0V/0XI7t4xmg6qXH3kD1F01OP
tI7tUTgJiWgeDNdhm+lXwI8TIYLpeWH8KGyyS91XkN5w2kT0k+DD/veNCSrK8XIR7HhtJaLGp4+h
BHY09ZAUB0PPuvGuv3KnBSTSMSA0PMxR8KUXpKWdAknrrNyyiFx8/samzGJkItIb3m373lNYss3M
yCE3HcY+Yit1ImKjFFHlAln8J7Oxbgz6jlHLB2KXV8leJF8afPY1s4QFPLULUVH5aVQwDZq3nuEk
xPRUHW7wpQ2syzUr3p7sK4+h55i/p+TSQhvnteymktAPhkkWX0kcD3RpX2oxomZbhRAKolhIn19G
O0pXNCuiIwbVOecgUMlt+NIom1B1Doieq77ai82CByAcKPIrN1x68H+b379yDj/Zu1jCnG6t5h5+
aMBw5si5xehI8s6k8nBqjjDBvdQkEtfLCPthyox4yyTAUIc96k9iR8TstlGz5e51qjJ78OdspuVy
VFbQWIR33+aPP+ujMj921K0e3rNp1R/v2KgJ0T0gRENSWJIPdd4fYXvid6GVXHWWLNu5MLbqLXfI
KWCX+s1pBOVnCGG13JiIZDFJXFMA7JjlLe4Ua9Huo9wm55XtF2fwMeNK0O/6ZHNZZCV2kW8iAv4h
ySYzMhJjkt6m8xWG7FDo+FzFfHxov9MlznK29gsHUDxIFJEwTZjVids1wh8SmzbzN7xZPRPzuKbS
lpDdgBVzbhgWSqr/N8u2VcwG4za9ET5eQ+i9Skmzviut1yddKd7H7Rhcm+7cZYBl5ZR7BZQqo4EZ
MXIv7xDCuz/d2SOLFbnSgKBLf3KqWeGf5OTIlO8+hXwYi8Z7IWFgZGYy56YfhWmVAlETqJ6BPSTC
vMYP+Hc4NW9zyWThR/RjTnaPxq/JAbuPpy1twRto0ackvfuDsGELCNd6PSGqogeWH1ra0xUB2Ggy
PjGsT7hXPdkLB0ekDvwClCkGexr0KVsy9eEfKnIUG3cpwy+v7hIEg0dTQT5qD82W4soPKIc1YsGl
pl5EXJcRQOyce7vD2CbdN3Za1QzPOoiJaqbg+F/ivnvBCRhzPbtCFpDG3PryMEO/h/7Svsj8xgfG
+O5keqny/zDKxI5MOv5/7KT10eCp4+g9obBSbjub/DVPs1pyQCiOc8IRt3lQdcg0vaWy9B1+S03j
w1ea0yIWpVL8ZwzG82XDSwz5Hl14IN5yTEm2zBlAMg9Ps7e1f/xQVUNEz1oG83A8rS4gikEEDuNm
LDEIS83mVtS61/lKiMru9LgG0kJBY92lGpdE+BqoxrnC/YpUmciNJTNfmtfZ+9of8RWcG7e5lHiw
omkDQ2naMeD708RqUhMktVyj9q9c1CW3h4+JZWiQxd/7QYW9JE9uC+nH9OluahfV5t4OzvOUpNDX
rVq66GEw+Clo2uxuhCEbuF0CBqIaGWC2CipGTUzuAlHbUn7ZPeCDZ+qk8xlsqrqOzW9F+wzvuASH
9XN8uZukRDwscdRjWSkQY9I4HXm01DWDd8Nk3Dup/vd4s8l3vLPBhBlw63cYR7Ayi0YNN7oEW5WS
mcHLWFOuJ39BTUj+m8dLPMT2Nyh4dGdzoxHiOv0eO1bLXRCIZjvNICVlKJI3KZsDuYAd21sqv2mB
vUW6fFw4USDI7LYhMj38x/enC2Lo7wqyLUdxKJtRzIYSsIUFtAPEW4LVj2nshUWFUS/cigPgKsaG
3FQK8ug4x2KXKHQT11bXS1ctEFsINvnKTl/Xrg4xUow1rW0FcY2I5aBUilBGC2dfjhfgleNiDFsn
aSzKw3edQALbRS4RxZcRn435iJ04rM1fWz9afgH9FUUKe+HKlBlmardGk4qodtVbTPnSmBASLQi1
4jEtCqq8KfkKZha9lwWOP/JNIuBseshKivb0gcLdcwSArZy//oVJ/+LTmjeLEmvAVkEdLZ3atsNT
7QhwmV+3ieZgBFKxn+B26g2bvqlV08uHc0wFDINOSSSO+/XDl8NSPHEvHFW3oo4JFStppPDS3xz8
hW5SBAFeTsYwgMlY6rOeTZtSHaVE6lws7daVLJLVCA2TUIgHqub7G+SOp4wPCzd5KeIrhgIAWMAa
f5q3Qct33F088coX0cN82TolnvuUZdW6Yoh2LgrVgNPx2//FE4TSTjswNFAbuggQroVrYkEUBSlw
XLj2WkWUG9RrEv6RYSAir8KoApeEEhrd94lw+4Lja8ujYxl6Z1Wta0yET9lzYyJmLowfdaDdaEm4
NVl+ROlrrJOZRszPuDE1B4shEsdqj7b+t5LwMZpX8yDAauaRrENpM0F//qfTsw4Ph4ToGOioT/de
RNCdT2tRBN/C9xtgz8d/wsRmzQEslUZAAOwy0Xp5XHeMhCx5n5WryAsq/EDbDMjArI+I/Fd72a+E
z9pE6opeytxFPhNsBGOsJt0Eb9O1uoLmrvDfXlrbCsARgO+46d66BJjc8PYbiPYpVCDsMtXuIy+M
jIpbbOfu5eaAtgyB+oJLG8pU8NWpyY12FPK6PAWeMZIWp1itE6gyFXS+8kL4V21Y3mX1orZK1T7t
LN9HUPrNyIccZFxq8gFyI43NXOnx88PrVomENxd4NmIh+OiTVG2zKcqaPNDNn1vvcdzDzfoIBl5l
SB869CUHf/HwAxh7osEl+mHv0MW0nVR6YUdx3jAe1K030KiAhM6bI1GWk1iKTb1IQ6BqrfMLGeZ1
M39qYjc6KyBXel+uQ/bvps+ZCBEvVEnWwitljx1sa/cr7rVN7OujnkDZ+TbHU3S3MPdcvhoC6uE5
dI7HGSg1hKOEJ0sXvrEEczerQSyqGk+IjCS8R4mbPj8AXMM+PVqrODM1/lFnY6Ool68WeKtip0SU
HefzQwqmfS6Hq/8S2FRQ1BQ+leiVv0Fbfi6WMAfQWCY2lFV/7qWHxcv2n8Ej6g2SoLpUTu91+SQh
Ipk6YU2/T/KmXqNTDPw/t6HD/DWRvXrLdcjLRQdqGS5Octn7VE7pCNOAWPXdwFMe5DvD/f/DJxcf
1WkNRvidBPV6OPt6guHBlnpoYYwQ0QE9qML77/edwOfg3Dip5yGuCy7LYaTYILq06qcTENL2xney
C5mOy31Ey6p4MjJVZ9w6E6jljC1EzDulU8nMr7G3//NJLkUQVlE1oiuXHg9F//xxUwKIZSc/fAlL
GcrX4DTKuL4TvbRzENmgsRxfBuXp0VavUdPP+n015obSp8ZxhLSjokFoKaBxrF0KLgxN27COdl8+
PgAoOP/we3d6jVa5Mv2soEce+QmbSZPvsp7UALQTU9DKMb+5gYXm0m4g6ugVkVZObdyjlzhRSxQB
b4rvdhFReKAxR2rxrRMTYbRa+lrDkvl7aru1tvELA4ha3p1jgO1b7ICBimccZ4hMqkpZf6Fst2if
J5IpVIXuC4eTVv20gxdJiNkiSgU7MkMZiA8OJvFrv3r/VXFLX41bmcll6HV5VVRRnI/2alq5bMXL
rxNG2m3qlMORymeMHH7y/35zJTyxKpYHxvO5z2AeAHyxI2v5frUr1CdVG3hE0BQdLCmyGuRHOC2d
VYrEMvEwCje4YoaWJ9qGI2LuaW03NY8IefVMhc5zkvC8zq8GUlRiY/uUZw9iepE4+0PZQ/Z68Ict
0Ff1m7tuMychhFZto99h7AOG08N2Ob4nJwpQQRh1J3KVZQMSJ/NdR7kBAaxfB01p/PnMEmQ86uLj
pSrQCfRG1WnDZ9CmxQVQ/yGBPHgeBKrClvZARLYhDo7DGqag+PzQQLsuk/S63gjmklnzRqCRsQap
syvqbFULDvLjEgxEEwOWwXMsE1I+e60VnPEw83Kl5lvRnyJJhuDjEGxA/0Hh99sNmcVuSg3Z9NTc
uPgonJLNy2dL4ZnSh0HTNX4bj/25X+jbWSOwch49UI84tgF4DNZQgF7/FVTEiXPYyXp3LecKWAYY
+3anO2H+5XVosULTXZRPmdWi9P2OrZgjKxj/4tudTeqo6aEy8hyp6pOABAYIVFWMQc6cRjdNfT9n
Ptr6nXrhQBkGTe6hyL9LQJd/2sVJ0l7Gc4L9+NoSvGN+tlY0a8gUbWadZU6wugwiaMzQMB3WA4H8
2U30JaoS5oPG2LmhOrNz8hHqPht6rwv8XcryTxJ+TcjVuoXQJjgjuBopvcCfGIvp/MTUapEJ0cGr
3M7r9RAS87UON3dmavdv2ovnA2EuPWXuGWr1mOy1+fa7bRe9S3gae12fYpBzs8LmB6c3+wREBzAT
SkjD4zEEyp8IdVGVab/bftcpbskYsUFlYsYdVkWCc2JdP06JvBJhO5h4ht94NtM7Usj1neUu7Yog
RxMjaHg/gdUsHCi2BlS/2e7niK53dp4uTy06TjB3LjrQ4KHx9dgNH9jtA7i94Hm8I/pydsi8VUEL
UWOJTrRD4sI6EZn9FpA3s1u4teiW9myW7IvB0xK7Vmnc/JTFrqbFupv/gBW+OD1DSd3pCsSqmiqZ
RuBizAqHfRLT7dF3m47BvcwbfA0OAChY7Ivbt6xcyFzsun70c6tBNnsCGxts1YwEbS9QVtlq7xeo
0BrIK/mi93SNN4UzhbgPbZafpFQ6DVrtFTDvm1vFJpNmzbAa2CVL/0lGlcZ8YB6LHBLLQVjJAx3g
yyysEegb/dS4AkQFdjmZY07l73j1f5YVwcFVD99E8XH+q1YE9ctG5xIWYupwz7lRsCNuv8qhx9un
A1WcKlED7tUcx04ugqataY15M1Q3+tgodiD4GHzMrGe5xQHg8PR6sTeDuKpbDQi+8igkFlnYWLYq
t0VSPKRV/dsP71Ran0bKkWM7VxH6WKzjYl/OcntNPi68cPvY/xGtf+x3zovKKjyKc8Wld4kMjOuv
pNqf+HQsEy9i5ltlPswWyOwbCm1dHaBff2NZYkTsC/YeQCZKmewIR5+OdVwS1UQs7W4P3+KBZ/Rw
oh/GpY/blJW1xzSM/wftGayIzeqGE58tE3vwgXZ7usLzTIumAx02N4ePu2cmPfmYu765iw69r8n9
5HJdpHp9OqLbRMsehhraGxP4Voo+v3Nf/gvNClgn+0vrQNfvnB95qr4qPNWMtVo83CALKATEc1mE
kkjuA5OzOerLs7r9yQ5Z5H/P7XubNrt9CerdclTQsPySdRyNLvXXzAFzMlKbDa2sgZBMYlkIiLNh
RoWvxyUgM658UrxyTvB3ft5wfDGEMkpCz1h9LxW693F6vtReewuv9tUJ2AOFFf+VGfB2tYgGxYLO
6mhf02C6t4j58QRB1jNWs4B8AFbHwsEVjI41OQWXIXK6/r2MLQI/b4Wi9NttMPhZi1j87GriX16N
LcPnQ5vnxF88kh/WnWTHqHCVctfzrWt/Lde/O+zSp3B3IHHgewp/qNrzUXLLHA20h5Ncbdrde4bf
DZliWDdrDpvwrYOPK7uCRTBky2eS+wkj8eKCJyeAJBy13v57rciKb3rmk3qDv7oBFYzdFjMa2juG
lpx/JHecSs9lWqqGjaRfc7tKpTt2ADW0R3bQ8fULPDBqFnZZU/rEZmdJi6wKDjCW0XhlFOoscEGM
bsf8VFlU2eUQIgkHcSYHo+K5G9JpbCFuSXbpBUb18uBgy4gErR/3cqfi9DbcOTUtwx45bvpZyP1q
/6PpGuN5fSPCEllqe0QGWKAOymvftaaaCWkBHT7JKcgS7OyDYWAPGJLmENIXTAm6CvjvobcjmSdR
0EQRRtV6wTaEzCZ7SWtrNCn+Papymlk4EJPrfh8cVQj4RHcVOZIliOpEVecZLkMOid/DF7sN+aAG
hjzu9InTN/0DpzrZxQRcN58xgFN/2twslm+/ur9LTv8QLRq4HoghgPRyOnSKldGOtxTCFe8thPxr
zYggktg3vAhjaFc/vk8aCyTDOVZX0FnJtzzgF7BC4g13e4Vfq/28p7pEycVlDcnc/hQ3XMnE3MSO
6/7BGtdYfKxG8zgZcdbKegQAzRwnqHGx1w74zfRl972O8HuU8O2ykWdD7svtn3oxK2ol5ehH6q5R
8xSsVk2n96iuFJXoPYVzRGNawTe/en/+oWA0OT6mrEKZocuwfYE8r8R4mHg6ZJN1YWfDtP7Y/2x5
oyAq5B2OX3d4zURaVRewd84Q1e6t2MCT+Te7ZzPctGUf/n5awU2GOwyDZB1SzSG7kTUqVqq0z5mW
FJ+lfykXMXF1Fmw90waZ70Cqe28atm29X7nZGTVbulbT/2IVtDWFLX8bk04dh12uNqsnV21y5EUl
hlXekvahfUaQMJnn+oiuySOlKUG/jqb1JlwyIivqIzF9UjxM981l9oSFjp5QxPVBvMbCHYH5T2Tr
xA9Zi9nyKY9J1yXZcWShb7co9IiwL2XF8kGVZbMr2lqVgjvIBhFuPipZSr9GDW0nLi9oyqmESKoP
e5n79dwrzbevfQLzHrQ+yp6f7G26PCF9kfvO9EHojXyb4gRZv16vsOeocc9o6bjteul37M49afC0
9wNwW6swucc0gvbaqHSWFD5VxTv/vfd/37/Z15g4TwPvT0gilQwpgovu8EbyNxNTuenZyW6OGk5v
8sIeslAvOdmVwl/hBRsB8fLnuswli5eSW5ZhZcplGLovleyjvQ9nt0nkjyV5joE7dWb8G4Qa4Nnl
ojjPG3DHp8AuqTgXe/0bwtMS8vwYG7AGjujS3ds91cB/jE7/nk1pwB5gBhaJstJpAKoigigBIrUl
53cJq7d2AnGA0YFJ7fZ7oUbFjMjzgPOVHWWpRJAt5A4yqCByZP56JG6t5cu7hOqgaDLne1VyiiyA
gyeutFBRbwZWEOyguDa267TnqZSuJta/KDVs2E2gvwNtg/RQTTl+Wl4aNAwGt9VuAN6u9lPweVVs
eK3emNH+kK64fRpblCShsAyxzxOR+bgji0aQ2fx7P6HGQG8iroNFXsVdRh6/Xg21n9/x7fgUB0uH
/lSSmmnqdy1exkBQXe5xHaW20L8p42SfduVyVmQWpQYMAgHEtXdCRnpKG/PItzeefwPzznm2OIEo
xf9c2/yOs4cdBk41+FHC1yC00mkq+wArRvLFzMzj2JKp7CYZXDO4en3EfgYw1WAz7/Pq7l5NMb17
Am8RzUMVFrgVGsrbnmqlQey2qiLsViDdvcOZ0NeLUgKiNK3e6f0HzOmJ64FXA05I1vqAU5zCZDhu
+HGi5+o3kr0SgVKQL6KeKzQhcwbTMsG4b1BswobDZMFmyv8+e0X5KjXvacngGybOCjLAOzVcXj5c
AaAI0x7IlTSqd+TU6T6FVsOAlKbxDwSG5GfF1TneMaT3++2Og7VMAhZ3SghQLyWpRv4ONDqSPzQ0
31jXmiHqRYEOBqi9bCHHhmRRpAQ0n8phv+UHNfeEgIyZ/0X5fhn21Jhu1Z2vKGio50DGgQkm5MyW
sIfefDA3v26C1hB+dM6QjieeROMmriSotPveZF7LweYdhK6g8ztIECOKiph8bIbszErg2FOWdeFf
ucoQfgTXYK9c2kyzicK8Rzb5pkBSt+ccbowV9immVLpVc6NjaJnX2JCKc9yCn/wzHhdn9qUvYeFv
iToxqWc02RdCu4pVuS1plUMNNql3pUf5jHS6sZctcZgxsK+qheZsdyOqnjQLdqOL8Zaa11QuQLlf
AQHv0kVUcjKxome/UwHV3thBn+DrLINdESBVE1jkX5KTfyymgjWfX5vbOeyjhjVhrVbZV1Jbjajq
H/vhufdLdHx6gdXaanuTb0STH/M7dZPbTZW2nQHOxK/yo8INGauvzgDvHZJPEkVF2iSZM7A3bDBS
uwU20S9KRs+BvAK1Wk38MO1Hf+LwtekMybxqvZhYe41+um6WAT6q9wVGOXj7noqrMGzqgtRbkdWz
rL+qVRq7txm4bZ+RuuG0HvYSFUo8SYBurgPZl489qLn/BVCAR9mzVETf6UHt9yonIJi2IEbtPjAJ
qawiI4CuhhkCxgauBPtrn/8SwodaLMTC+ARPuhWWOWLvdeK/si8GT+7kJGbmn72Uxkr8H80Q616H
LGxVyYVqHsXkwCJ7nCHlUzwde5U4kWwMskw9WcI4ktl5FyQJJXQCKGhpnvi4k/2xeW8Cg4lpr35D
gUsaNLqx5nuLXBaNGRtE4pvl6b2ln5tUPl/zlha2Lp3cRAOlF2fl4oLFJ+jccskc6VPtu0aGCNj3
NHDKbDznWFvIMP0FX0Fld9oWMp6AE+MiCSF88OdvQ5X7Fg1Ftq0GaBnkkr0Y8HUODBISAsiJHa/8
3O8mZnybqxR4TnQ+ULnHrBDOt/4d8uTRe1X1Z7ijQ5/6tb+RlMc5SMWKR/FRgjTYNvx4xbbFIXiu
q46r2EaRixnCZqX2dpklHXjlSZ2o6zgkJ+qrZslP3IRmkGE6GdjguYfzIF8NcMANK2FhTza+0SMU
nYFSgtDNSuT8/fFXUcimj6DVo2gRmtzUg0JxrTYwM0PSe6QdENBTWMnIpFGLkRrUDxK+mOH5SBu3
UA925KrpLiQBOK8pKW+//tRCTeOF/M5XS3l9yb4xQ6o388whEX4/i2Fp1QNdcU6159Yu6uwv4vCA
+ehTTc7/MpyB+Be5kcA7PD8u8ibPGc9bvrlJk2k/TwnPrarsTZXA7gtypq3Rdh3Y/BPYtBiyKsPU
rRT80G5pUN6puExN+v0YrqEdz7sGnGunAmrKc76geEaVjhTPq5uvd9uNEZaveiZEt7nyTdltTwun
GjVRqvBbIk8MlYKmrJVPET2Fgsk4+cedhCde+3s3EYWbmmXXx5eCD5rFCBnyqe9IZx6LZadGb5sZ
TiNc3xyAkXfFO0UtD5ghbl+6dp/4rIcTprzszXnef0rGs8TQmt03/RMD82CgbfQV5hSitYXP9qze
9ADENwHKV0o7SOGD0sPiLpe0LzH38tcLC+02lhpmW1r+4wHwOVXIfpjYakexdlLTY75NdWcJfgnV
Q0JX+LVA6YyeN9WdDwmcMzqbo3khIroGEYURpTwtOvZdCfnGw/38clgt+t3hzid7gmBZuDO2MIQH
Frz/n7u4H1ZdRCIIqPWXRltiio0rJWeMrxm0nN7F8VsDmsexR6TGMSmLys+AISC0Sn933GxE1d/J
NN09axCQTFbHUtwbh/xmpsXLMds+S5cVIthMMpvLICNWmRiBHkJO36fuot8QDFg056C+XfiiO707
4mVdPlg7PiGGX6HVP812DsYhAwCayXlrX0Z54zT5Dfi8xJ08F4wTH3ZMwSe1Xc1o16Edurck4uLB
qLaXdNVjiy+KNH4pa6JntpCoi7qEejSmIHD+bApF41afL902T7h4C8reI0mVL/M6nljOBhaLDpjI
5qkSJVo1ZZ8TC1xfJ4Yt+yjXjNldrifZJs6cia6glrKcnm993SqSU4KFgVU+tgEgp6e5Sl2ofQ1C
jySGBGsioGqrJBYh9QIFdVprKGN4bdcU9JFnfCGK88mA4dThFqgfnVkjHrzIHPobUKS6Pu8BQ7Eq
vpdaC9ee5dMSyFAfkf1agQLn4Rbrsq5G3qwZ7M16ILPiv44r2riTXpBU9reDUHuDvPFCzR+p1982
QLBCO8XVMoPVL4qmQlARrltj4yKLQwWNft+/8WW1w58xSqR9BqnUiqZn/j64kyYsfr16HIgxADEt
7q047fFjmT9XAx7UpyfR+htZ6GEdxDnyWbC3ldIVXV7cUWOS634UG90dipcTclOnw1Jqhm7kHrMk
nhl9epLCtGWeVu9znj6BDL2+4iwoOSX9b/VC6pmtNiwZ8muebpOhqy82nPWxRubAwshQCYOYz0TZ
zCthbAPnjwJffjbFeBxH0rfdhLzwijAfic9fHQ6+wLWESf0woIjrCdcxlu3yMyXQFjzo2SQ0ao8I
LP5TozxhgVsRpikRwECvY4+X+botjb/Nl0+kQY1TmNs4RdQ3WNsHM9W5iVvg0rLhaBsmaqRfVsmN
QrbqGj+qN/smvXwWwthvmDEQvHJZFcauxqLlnZhn1N/9Af8jn2yPWGIRDfGcnlOnH8hFuZkg+s1h
cIjpvDsUZF4RehL8qqAA7CtMOocqFnx+6G26ifknJaF4NMEGb0IyZfI3gXqRaSRhn2vfFkwN0GvL
PcPQgfLqPuJI2FJco/rbrCfSg3gffdr67Mvz4cXUve78UMgi6nIcPym3gh53h1U7LJtm5G3OMmAq
+Xf7hkNWr18tG9mtXeESlljlGYnGwwtpF7oBRuRZKx4a03M56mJbdlRHi2V+lD3m8veKxC5l4vgw
FIlyoaCJWS/53gufU1lMgu9uBjACb1JkbbHfI/wwQyMvx4xRKdwHA66/euZGZxIqOsNfdM/zAHQv
BRv3weuggWCVxl7SbiqOhjw2VkYKIdK2Snr8cR2jnZin7AbDMs24QV2RZK+jO++C+/dto8MPkch9
eqHcCiDYM4hrnx08kEeLWt0nr0cyqQrewlodQeVRmV+mTQcTbW98ypY/wb9aVh+9hh9TuMzZ5psI
MyqPx7hABqZJwDAeRqSQsUKlWeqXVmpGRvE6iuM0t6cy6/yWf4mTH7R41dLOoPxXMkoaY7zJPzNM
uwMwn3llIM+xd5aFz2wuVFq956+LGygRsCL7f2AJT7XFZVB97ARiSMBgDgwuiCX9ltorFZgkgVng
IDX9Sncm2xEhsUanph32DC5KrMTKfjseV1dCdGCOs+Dcva/L+zac2v2W9OBNWSDtvbB/T2886Jey
tGP5a4uF5mMuopo3Ww1EK43zSio+401d9yOgqpazgDqRkTpLTJDjBDFBIPSrdcIhSy34Pdnrcq39
tvoBSvVvnH9QlXSiXL1spnCrfwV5ekN2Fi35NuBS6NOEzpeQ8IZfy28Nu4zL8A+hkv0BbasXq6wM
txL1inIe1gmkG+OKKaxgYZgMXvO6oOVnDjty+0U9U+jjmnO8hihNnhY/90ikrQxBkOeXbpYsxyx1
MdY6zHRE4ToVjHi4Q8SQQL0SuBXVLZTw4zEcfM5YFuSy3KueyA35qc5N5jbmvYzMcHcvpaa4GP15
bg0ar3PFw717Rm7upuPYkv6Zkyc6DGh+fFJ3qSk5UX6caEhuaeVojCR1ROq0k+1/yvb3uMwExoMj
q7/4OjEMG1qaE1k0Dn5vlwI8Ion8r3jgHtxuzzfBadNLiX1WiLciZ9dxWqB0ZmEclvzKCJryj3oY
4kuaYD1qLKbLUvefypE0gcXVrSE2GN3l2Do0ktKnwQpqIqxz4DQe+1HuJ4o+vorgKkLYRNgxrA3m
8L6gPZ9qe7eFOahYHP4hl+tmhdlK6b67c4fhs8/rWQqwvobTpUr9uZz9zvwIef3Qwln6O8UjmdiF
Zy0LRc44cn7l9Quuxcn3J69psj+psuQimdr7hd995cfkcfdWR6SgZcoHn8U+dM6f4WbG9fazcr6n
0Lts9tG1Zv9rN3j05QGl12NKSwBTZOZUyXPno/O8xqTpptIrk5uhgW0ivcE+7DeYWe+7C5GR59xm
5MhEEnhI33GrQSiPp46AoI+mymmsAQA1rXz1QLDoJdb74ZQEstyC69PyeDsHJAvBfGe77XFcbAaC
JOZ5p00wxnqeZh7iVL3oyM720t5bf/xetn+ZKVx5djKuk55cVlJvn6Mvm1n5fBRSQvB0u6Yu0bV2
xzO1MKSZQ6a/ykOQUG30twwL7rtfxOWjgQuk+lIXdrDfcOXelAFHKB3tAUxbEFSkfPl0J6BkRMDF
4i+rr1sEvBVvXCjlG3NSHoo+hkDx0b4DNF52ofgyW3vzIpS/a4+KTZ/fxKupwxiHfa9t18SOoGNR
qgAdpbA80FLaXz9cGMDZq8kazxj1WALUUOOrFCYAl/8kkWjLGsWIecQH4E5aNIsA4kp5gBsHFceD
e7f01J4NkjXuRRuZs+roaVp0Nh57VtJxKqYtGTPJGBUzOIry9ecjfBxSfJ+KhFD3O90EKuXEVTIe
YJJ5xVeI6Zj2mY+wQNaf/yp+C5RrT8GoT/DbamGJrJ8wPBBKdzU+cezGVxCjq7jBa92CYMqKWEUp
s7S2fNJ4alZsunmMSsuRaNE=
`protect end_protected
