// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:49 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JIGKxwEfDxaHahqJrV+aRdbaGyAZJRHVV6ZqvEcCvy9iVpa17oBcf2sjN+eRt3qB
r+S8z3H8Ws7BS44ygeNq4zVf7SX8eC4DbQTzOqRHJHkd4Ir6tPMSF+aw/ugyFIFq
ulAMcdyFFAYQ5H8P+naSGuVgGUb0imxFki3XHYkYiGU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10720)
ALgaVpggd7ribGz6xnvFKCsNoMGeBfyUUoMR2JlOR+/6DPooC6/M4ic7Zg7eBgNX
1axELPXmjz6ezdsVN4lD1gWV23hFnAmRYytJttdLGevP9s47bWe5aysprxjzRL9V
XWnuF41ZXq2c3FaKRoQ1unNo7v8mC+cTvfsxXiNxos61Dc8s2UYqO/t6LXIoSu/U
bkDFlCyJEIeMR6zf6UMLqwjyr3s2D6LDPlwebnaSTF/sDmt77+KEvJtoXyVQjJSd
V61uCFFByQ7+5FWBdJ7ozFow5WNZG7AhjkUACeLz4kcxy8ryx+GdZEDSoEL5AytX
XwNn/ySs5a44DdoX/UgTANvZ3mcIHpqCTzIA8iY7MSEbuSXFQxoClR9UxlaNNPZa
V+ai3cE5WcLQiBmaESquNk0X+zFShERdnxNm2NnaLh3Z+ZpgBQKsSvu+gLjVVyAg
4aNbuSZsHGaVTAKcGvPbGOMzflDMEIfq4HRI7Tp1izZFZUGmMcZE5NHgKROOjn4F
vCmpuyMW0kFke7gRt9FM3fH9mno1Lv8iUam0V9zNd53+XhZXE1XHd3oTj6P0X8Wy
WlbuLsjPgrpfsFUvWjUmht7yqnktfDVAeJJPpyMnj6jkJj4kfLy1a7fu0Yoh4EJz
7jK7rzZwHJvEkfBLBEh4skqEvFGdMTntZHwKw0hC6nhT0WhCHoun0XW/vTlakISC
CTtxgj/Vo4XoIDe8JWwVjTIToBMgIIJZyaLH4ddhXK0U7nzniN0nEtoZkjMeue21
ADEY3I38m1DdFpZVuxTDWGi4slIwSR3RXVp/p3XibYfjdXfwcc1DsxRMDjmOBKsh
QiRpbvO3F3/Z98frPZlwzbgbpQba71Pfl53/kKM0JBsphNuK6QkjrDkRYmrBq4Wh
RHrovmu7VD7ks3eRHHZii0CVRZFBfnPCBDHEzw9vjCdf8jZ7Z5g+FGcYaUkf07ml
2HZsL7uQ53TSQnzB5m2G1QuVkTWAfkhuVEyghUygT+QLN6ZBkXcFFZy0eS2kWP0R
F9xOkT8PD9FvtTnZRkz18w+UwQMhFTNy7JT3VVAMxaZ82S/folRWTRGeshhfqoHe
Q3qbk02viQH3VRpSAXTsQrCEbdbGJAmSHBTntRleX6cjtsois/Gw5NiaWMTmjQ1W
mlrVRuxHRIZVYrMLSxo0nqAmJC9AdEd8BMlCasviRITFi8khrlRdS+IYbDNTVCSQ
3Y/0+BNlJ6ZdoFkBp39fUEkdZaqA1CrKS9Z046/HTtewnhXCI6kprIS2Fa65Fl3R
/Z5CMhaHx3XTkOa42+Q6kSX1vhlbbOjD312bjfkDL3iFXUwlWej/x7CAHrLBsceH
nJoxchL3xXyH9jdksOel8qtxcxMQQJYSEZPN7Nhz86HatwGEZizreLDfdcQ2M5go
baUT4vAdfvwFj0t4oc2cOBggQuFHbqLa55iMZVDu5H2OxCfv0htWVCYKoQTplDSx
vpQuFah9eVxiV9gZAfDjOOAX+7gJhokHxJY9q3jizl+DUjX8XiH6f5U3ew5TIaqK
3SXzNOCXpmFz2mOHZwGKn0n5z8rQJW+QcH48NyX+cFY5QtNorzCi/+O3ZkFoi+uH
p4ADf8Q7lykmAvout886AGghI1l728kyrXoPkj2VAuTzf2MTCR2+A7Df5i4csgkS
W7/5h5uP/UzwuGBJNC7g7Dz/axMgDPFh6BP6YmLkjl5GV1kvhSMOXeEmGYnIIm7Q
OpeSksrmgr17Yy7q1Hp1u2VOD6aCzZLbRmBXVRt46tsKDD95ZJZ136JvMVtSGtW6
mEIhFg9fRXPT3t+YHCVpX9f9tq2W+l90MgTvps/yZiTnxfrdjgXy/Plh2zfM/TcX
+1Y+gkv5rOcvlof60A3Q4/rZK6V9RflvKqBdQJfbZkuQaFTIl2HHIMHJqbk7UQ+v
4ju0ru6wkGoRWjhmRSeVbUHD/O1oGHQ/71sXfQnxqJ00MmGiokXWbVqnGAciQLd7
ReILcTc9uq8GfJo4nqvvVd0RCKAIKqaobyTkoBZk819TtI78oQHNz3n1sFmz1SFk
xL2WIcwLQbhoEdQ+LdmqWbxbJWOMBWfrUg+fEVm3TZnp7QzSqwqm2Q93Rz+uNSRP
7LPcFhM+Fe9vi37tE94FXkJJE1QzR39VEc8LwFEca/ZsLaCnyiEdPCkgtN+6OwMc
mYhC2PYvCW64NaWbi7vguBIlnSnCoZzD5Hr4Iuo8YkLOOfEO6cYOVVEIclVdhFEU
gnAh8zVCYwU60xaOCAPly70JUUsoMBJi48GqkyALbfyMI8YFziW90091fIKo8vo5
ThsDzL3TWv2zLZxeuSPDs4X6gLQa8QQ9ljZEIz8DTRvrAbyVuMRxNZmeQWn1iwgp
BM+Sqa5kq13h21G8ieW1H8kaH5WITSh7yHYyK3j6qXZ3Z2qsTzmeeQfzYBtHn++K
zbIZ2LaqudDw94ATkcXppIOiHrOGIUOJKGQIfZowncRz9QWLXpDBZ8262yxRY6/A
K/DlaCDsnimNg/sWYOOoS1Qdep+1HZm43e3APj0CwEvKFxq+D+PGYMwl017/mTkd
fh3pPHw4PS2Oz/GzwwRrOPQaYDDi+GwCeXvolPgYONQB6Eq8kTfc6z+5s5/HjLYB
vz4gIwxoUux6G6GGJmAlQpWHNl2JaaakcPzEBkP7AI3mE1nBUlQ/RYIPp9CAVUUs
Q6YaUCyTRrqe5CUj2g0GYIpoDvrv94BdWAJojHJOe1NtLWMIehIkGw6cJlDSBhUb
aIo6W97QHjFKn7dh5BQLKShmjlGzlPg6KwrnxbKV+HTGT4TKoBr7ER8pB27EXHZi
B/5dudLGSV20BwHPTHtNeAfSOuuXSnubUvN5vq4MDrH/NIlORBox7ftapYsagwQw
tAgJyXfwkWE4xXCm6HifCrt9Zp1ZktoODPLPEO93H4+Pjx22e1DdefnJVwlKj0Cr
8tMvX0gpjmQob3ak2Iv1CI324E5HrSMbAANtJk6i2xJ2QS0b7o664AWcIcxInLFz
A7Ccu1nm9/kfxUV3nqBwBWF9UyqeGunS5JMrtY0+Opni7t4kSnMQV/EDdx9ktsA+
uUZ4S+eSFgnM2AXXO77wv6LA5NbpNzV7pFHzDyEXs2vsXSj5koUWeO99VGsmWCm5
/cZAohb/JHil2mVIMksHU8gGxROyXLhvQIqvkakMwXNPLRCMhTvzjNjPx2kZcook
h2mjXm+LAri6/NgTT/RrB/dAQvji2WYG7Y+WKEVtBnThwhTJbIFNacSsciVrun4+
o9/lojKEUx4cvD7HekDBKs5CfNRnc3BORRBbIrT9bjcmW3JnmgFZZOutHDdK8Esv
hm4EvQGYvDMW2HiJoPPGjtYrLZes2HzamTWRf2cN4RLK+Z66fRlRBEsHG7LSZymK
wbqWtKlVwkUNxVTIWCM1mDbpA5dmc+uT45aV1XOREMrlBdwWPnPGbalRffJA9RCp
BfHhdLWP/usuc4Ffnc256GHe08UZQqoG39q7e+wJNuOWTOESixwfwZNxLyUX0mhJ
YffaymxsSovl3HR+aV87dYsPnx2YbokI7mSkL+5x4RtXk/tzHJdQu5L7wOdgQrwv
LfJuw4VnT839W+yjRBsR8PuiRMX6q7FsZaIP9oIxzvtXPGiref2LkCabBHsds8GM
6wbTT3ZionMIAOsA/YYlOX5r6578oCqlZF6ATk5DcfHVyBngbz0SKDrwr5u0OqRA
6auKXxyHl1/RKGqxwCa5Jjyj8HPN0HY3mwjUswFrvfxspduw6yvQgovavKU0u33r
Aoha0dvYKnm25FeiUYEx4f4b/lh3RqV9Mgko54+BbYyMNoeyRMEHsEUXxz5uR6gQ
cRoJPJspuDuXZuTy7H/iml7ciCIVooiQrCNTKanK4EuzCM+LOni5UqCxpbrEbaeL
hF23uQvIliOQ8uCXVepCN0xu8JF5Rlngdh+IL+PtOxFIJ9QeLsx4e4ZiILqO6+HT
fdJw+spxeZyus1LIcjSQOgdghQAtQMZkXL5iNfKnKEYpA/27uO4HOhg/D8T5Fu5f
Ngv6p+SgkNXN5ftVJ8gJuOzDZLMLqxesrZag0+AN4N40d7dwcTaMoBFt9GV4We04
pkg2MatGoEhxjIoBz0AI6P7TessTvFfbupN5WB0LJEu5bG897zWatPEeQzRxcMg7
QzWH7p4IyRjmAp0BzhDS+ECTaflnU6zLu+3Jew0Fy0F2uLUglc+0tkKmXgFyQxvA
Vg85P8diT5d4Rn4Z5Q0c2Jny93xhWx9HKIsBNBy3ZKQhLhESFZMURi00CXTOCBcg
M2CUnmF9QBZ1xGtXILyVbBg66CSi2yO31g6lcIcE7jWzCRVRhcvSkLhsBkzOe9VQ
SXJxL2utBHhWYCfO1WTjkgIR/9GYmuG9tmheszFvUNbKHXWE2dr9EdrpuEf2rvcn
yjxWjo1MscOoXLvHPulPBXMb1JfnlW1g7biWQTUNxPUrP4VcD3S3+Jg2es0dYP9q
umjOn52yzXdEmwPgldGGBGzkQ/FU8D2j9dT12VOmQd35BT8nRuP6e6JFewOHPjpB
+OIG/UVwo1YXui/v+dB57CQBvcpNTwZeuuVsZHhV+eO++q1d9ty9WobZ5k+vEhr2
Ufd3nLiUIuMvNT12fIPVx9dHa68v78uKpVBLFg7GhI7IFRboBNBN7jzmWy/t40gy
XvBVtUJX2na9HGQ7+Nx1LrdsYyrgUCNdkztrjn03SHYiiJJcJN/fcEvOaylZFonj
iWmtrUW328j3INktbhkKZhkMtRaQ/+5LS1QUQB++7iB7Bef2iTSjbVzycpZNu8Cp
LW/WGuoPCnpALm2WxDQAKYnFNI/EqtoO9yV3Mvrq1fXuMbjotZpk3ahTknq/Rkkb
rW2uxXHM7kJZH/c/TmuvS2Q4EN8NuyWZ9c6/kAtjc8gy9BQJUo7KHsp2n4G9M2SS
/9dO9vfhOhBli+qZfJUuZxLUl2StCAcQdvoSZU+fWDGTw//3hTKZtXo+Rp7ROJoC
bCmpGOdbUXe3UAoMo2Umi4l+3951my541U6mjREGirtlxNW+vFAveTlRUOrpthkf
J9twYJwXC4ucH6RUt1prFtgejXR+CJCKyTnL/F51CmoLmpzMpKa+KtHSSgjWvffd
ACa7Wy1JslviCjdVhiHOiEzDQzUqGHJpfCl7+wUUlTplymHXOvImga5H3srd4WWB
ozmeLZ/z48yJsFEUlYZZ2RKzHab5poBfXGhvFSvGpjM0WuApteQSHnsaOHTAZxBL
tykHs2f5hPpmhILq61B3UK6lfj3lDEQsCywQ440PF53azF+63E5LJRKwYRj3Zv3i
hcIXICzYJru44Xh+ckC3x045UF+tLIr4gH70efRo+HmeBZ8HYejMK3GAkqsOAcfL
E3/jw9saHXm56AVozIWhq4CuonBXEOlso/cPfmsOTW/Y1iEyTrMicDtHU15cxKUt
+IASpzh98DpBmECDMUZKWgVWkxsB29JjERQknFlBUDDwGnD9me115E8m37/IEGJd
Jok3mXshD2deTcZUNM+ZhcMyYiObrWccxxsuTPppC9UhbLsicEmCozDXJ7mVSjv4
U7OcEpato1BoJlxIuIwTLGGVT0X4t6kd8t4myH3dAc39zuXTXRmWnX5Wzs8Lswi5
FTWxieTG476io+Hq+nq69DolTv/UbCHfH1ibA2tvMEUlcvMuc21sGBxBSpYzLiIO
sB8Ub8ZLUK0mzwWK81M9lX2+oR6/UxBLO9d4q2xWXLV4YnXO3H7SRmbaz5VvoDDg
F5ylBmnCea7Qy1yHb6UqUepnRT8KyImBFi8dgiLRiN5QMW30JxelxiRiy1g/Fu4K
n87Yb/8Vh60LM7mZSx96gHdodUvnJhdg7rbgMqAgo9lix4kh1FIXf6YdN0cULYZL
ocHUf4E/7GhJYZ/vCZlTKFgpgk2TB6IDkT+1amcpiZCkcBbb/p/KtOKcBPNpTqZo
xC5u3EjZkzMJ9CwBOebu8yeWHRMY0iXZa+dpKrSZ5qgDC2MtbBO5n3snp6OqaDoj
oI7Jz44hdhkQDzJnlpk190+/cPmnAK/LNfoQLmag8uZR1jjjMlHbTRzCTdpnJjdD
HMZxSdGkd6dJOVGFGML3FredetosRydBUIDdUpBqrKyWK0cugCoEcyIX7LN6X9GL
zt1sbrO3kQKXII2toksOOKndXs2QKKL4bt3zgQmUDmy0lpABUhg2Ijd1jNGoLX2k
B+z/iK9oLWz7USQnCEhgDn46l0itN+gfR7gLyn7qVz8QdVYUd0S7Ksp6FoC6X5wn
VCU71ZJ4M0HkDXOn/fr8dk0BYZgB9Q2ow23h/ywOVcVSeijPRO15kH3fo3j0htBk
Vx3r3SUJZd1CcGUagvDnccImfSrTsXCCayXqZq42S2UW32H/Xt/wjqpVxZ0D1m5a
fBZVPayoeu9TnqH9FpCC8fH1AhhoCWjH8fPiAjY0KXm965rIkDC1lhpHZzYIlpHZ
GeypOJ3HQrn9xkZ/6cmxgaefbEQZlT/B++1q9pyl74S2IyhGsC+m4LNndOajisDJ
li+AKXaJxs5D88/eH9E0x5KHe5i915C8xTmjNW1aXR3CSk4/kFXqXnoErngLYPyr
gz8Gj+tBh7UNLVW/hPjQrIrLnSAzM4EpRbc1VQ5lT7BKsiYiqWNszfBf0/9uihCd
A3lDu3CKPk2DbTKg+4qsmik7AncBPmL9Q1En956vHWkzJPwv81n1Ofv3aqft5SPE
pbCS2WVPgNxgz0NjeDb9OyWkZezZCVZngmKY5Ttkgdf68S+r/2XttUgGXEGM4IA1
VQxaNqJeJzJUTC3ivvDqm84mBTMKuB1BK2ol6k3LhIj5AmtaR+oUf3ZQr4UI9TxY
hrVc2RXQFTrgS8pnzVdQnFBVnVGNEHbTzoEoOjLkWYMqPgTQo/ZBDXbtACThqTIS
B4aeEC/9hkWH5xc+1l/9D1CjRdJ0pLJpZDnahAjinTLGJ6zP5qwvXBAf8porS2du
sY67XQ73n2zu1hfFSZF1g+CrIeOX6/qyOVLu346PJyIvvJSJtOGztO2ECjmLHefC
gxl8MVpZgs2lBqsk/NIBDfzFKFExyxXcmUQ8gxfH66l9Wm+DMoIRDAGWtex5bz0F
qgOJuC6JTexFP9AqZ6sv28HPyw1jI/b609vrmWuIj8PcNk8Nmx+GLaSYxF8g4jEr
E/30uVzBmemEKRdka3koukVkSkpprqPUj0yAmeXUYtXQXtLFdBS1LUTBWV27E991
wb20tDlccBbBW6OFAQTlz0jXoM3h65uTGkIJ5GfBktuJ5Z7zp1PCk/zGPhMNq4T0
TtUTAb89QjnITr8WCTOMBWLECZTm4SEg0h/a5ugp3sgcOECPTpXbU72jsbN0t0q4
qmWGgMIUFgXzWzXN8ICoxhjnApYbj8knn/DzqKqXhRa+5cOXhYghOD2OCWg0Xw93
RXvRmEgCrprFcRy44EVUyAkXo0nBOJnJajEIu9nFUh2s2xyCHrYxfTL+RZSA4C6U
doruAXYDb/fISVBgFmSvgp/ffknvDtDlRO5fj47CEyTqony1zocQgc6D5IkIEe2r
i8qB6nkuKuzcU/HLRMvBCNy2IUk4oVg81fowrS0LkvWvOBTfP5er8mSOUsts0WE5
uNBe1Lsmf759C00ztp9j8sybrBr8GbBE8u3xsVFzR8iPTolnPyFxR7MNbsohJYQO
9RQBdTRBa1NjMQ3Z88BWSaHSvaNaOIw2y7Y4akuXp7ZpAYypVZs1yAPtGNwBJbnZ
olVeb/duJs7jVFlhEneonUMYUsC0pOb86iHzo+vc1UAJzO9x9Q0FHyO81TnqmGz8
N1KL5III+tKD+JLiURp1eS+MhTy7i0xHFUElBmpB8NVVNRQ8rjipdsNVEmfmX4s+
BHW7vI6GYG3TOaixlbiAS+87iRa6P74BsIvVEhOn65KlZPfBbcBeIhxba6lc8qT/
jb5+PcmSFUP2oXHSOeLRSbcYOFdgPJiBJFFa2KG49JLX5v6/GLULjQcNmSbylbTL
nmQ7aPyN89wSjDcMHX62XDzSlxzu0IXTOu4rG1Jv20xCZnPOK3Bc7HD9RiF18jjY
qJHwFLDG/ke76zek2rSl2OyIc2+sxjvw+umaqoG9BL6S3caRA+hE/odW+1WjEG+w
svz1BIyk9kSSIzx4ScysGidX4aHGpggjJPkPLS5TM1lPhawEYveR3iicLoxDAi8w
BCig+va2EioYghBoipVqfqAp3ZZm4zwEvyM4Wgr2CqtnynBcQsEo2qMT98RSaa74
ycuSqZr1WnvU7GraKrLZdnjvlGLVuDpMAoX7an/4ywQX9sFDrTtLnqRMVHEgAXQU
+u7urQJYdBCPtsL1pp89/sWEYjbkPNOCFoOzxd7fzpPXNrrOT4Jq8AGLTz1uzzJO
tsUb4bB+zVFvUeh8401GzZjqmczpCrQJJxoVvAqclVc5hMBYuYz13iiUUQoCsE1Q
adhAQjJtV4cY2yqIYbJ5U7ma/IrjcHCcvEhv0qT0vq0z2xWRUqCoSrmTqhJq0s12
QndsKKn3JW4EIvvI3jFlOJ83uxJiyD7PsFmbv6Fr0CRL5rn5czEYMhUPY0tuAR7R
Rdu5Pb4FUMrl7EOoH0VGqgotSxGWV0yo/r6G83Kr4MkLpv2iT9U0S9zJtSZMiaFj
FoZujq574BzjlEUCP09MwUK0w1kh+B3M6ijJ6XxJ3UOtvWyeo3U8vEu/9SMPBJv6
1HsTpJB6lRGyu8NbMBxybbMxmT02f8PZky+F7NVZiWosh3YfxdGO4TvkhLmESXXu
skGyJxTyu1lficKn+H7MHjliHLnpjZeYgx5nfURUnssIYPYekcG8VeqiVsMd13M2
jyasv4JnT60fPdx3NbSSIBB0nyhBg2othWKw5nO5i4Z41pbg9X7DZeLfTp7kjUA/
GPqc9g7KXT99n4O7iUnSnMsX3597YWmCwMPtI+C1DBZ7vc5X29MRy6TOBUq9s8wL
b6Js5S7QT5nkm7WGjNiHRru6ki1q63jcPJ6xhR8paTN5mXf+Rd75NRHaYxcvRBh7
zGYVOpt5GNPOF8qJ7XGyNLhY56ctSNdJ3eaBKapvBavbYknSzX2vmLAWDkaUH40/
QPUq1e/OnWCIa46qQdb+5s8c5Ob5GchURaeLBkShq46ntZPAiDQS0AUXISCmxJh1
pp+aFAevf/QA5ewMuqnsn7J8joJhcQhTOsxwKf85II1Ao7EVTBb2Z7XJ71r4Vdkt
NqOA28u3qRU9U90cWSkSu0CNETPs+HjkpXukKTz2d/3aPIKEcYQP2+tfXMA4jJpE
1d2GPHObnA+rc2lRsdkJi2sM8/xuAcOIrSihZA/Ptg8q++BEZtBDLgtLaaD3+QgO
2XOfkcYqZALi4y35a/SyVQ947C2LOfDdymAY2esFt8sCR5p9qbkwbdkHJrjpgUuj
EwFsxsjsYuuuwC7E97oLr6bKHlYROzkACGr9wPFNGudaDzhyleM+HnmOi6YKQE91
HGFSMJLSDL6pPw7AV3eywwyV4xzA6Sud5PLbaYgXRneVW2RvQXYPzIhiyPhGKmqV
A1wIzVpkA9PRMQR9nO7LVKdmNg1EY9M+mJx68URZRQMT5XlNqyM/ZEm7D4HS9FA6
fZf85fe23FIb3CwLdRPFALJCFe/yDjoy2qq7vfN5BKNT3erULbQtogg9ttUkxQIO
Yemw6VEfP/s5YwXWukRgXLSlFtZL6y7Bu6hTSoutfhctZz3875HiZmtMcq3wy5QU
zi+EKQCcjXPAkw5NX4Vww3GMf+AuFns//3XBl3NI8nz1d+3wWcW6oj3h+LJDJ8/Y
yYU48psae81ddvu/fejSwqFydYVUCiys9mlPcEhO4RzOmm5TlFua/RRbC4Nc3Wer
cKnfTJe2HRg/BaTG3PTbBl0oqs8VhyGoxvzPBUox8uFI3tMIqN3AWOv5vYSDGHkR
8G+CTC76xBb7oun0/rDzdesonksC/SucbhvXEu03QHzwRjtlvQuu4TsEHc0BiQL2
fYQgtGho8rU4/PGDElF6ODfES8LZSsObeAvyxR97f5a/KkAGd/XBc6NEvd/p72Xa
PBCcnsiRtpzlBLCkztoYvcnnTgFcRF6vxf2kocZXAwX6ukciqpNcWuvA6kcX129w
cxgkg9+accc5FDSNMd5sf+acDIrnpgRLZRrIY/IDEyrcSfd2S1UPDH8PfRJCsnlA
EwYdIClqwYl6tzOLLk+FQ5lFyJKjCVFeC7W4nX8g+rIYEXcj85l4Naqcvb9k4MVT
BjReGKbH4fCuLaZoDReODN9pfq5z2xkMS1uULrokuO23+zBiXHpJevPXwu4KhW20
pU6W4Dc2/vmzPM+y+GkjtakPolDwzbd1UfH5voEkSXcJsYPdm1WvAwwVBBGqz32F
SwKWbJtjiMTKcsZ9uO3N8g19Lo6DOgJJnmkF4n1s6lkMZEcHnGMwN9czTinQJyax
7AWf/yLZPXjo95ZMLH/BCpq23s9icpt73jHwaKEpRVto0bskFyTLUTniQxPcg7Z+
2uShlNdfls2BaSQEA0xTzcN7KvkVGjyOm1mbJOwRL7yFUO/WRVQzb3mNQirbate9
HhSOnKlor/O4y2UKd2sEPSTU1zEE/IdA43RCO5iYXSR+r4/JHfO2m1t2OhK4Q42B
8ZcqKaKIQupHcj+buNUeAUGPSJ+/hWKHwxXaeODP+0BpXtMPQYwq7UNfBRIyvHsi
nsnEksD6j5E9ylnszcbu9aVvIVcbFrkbrzDCNEwU409TQE2iL8HB/qBXJMtg0rj9
pfeh2Sgl8IiqKJ6PvaOyZUo++p0lcGPkffpDtDzdGo7Zf6LoP50yd/Y96YQgbWzx
JZcc+lV5a364FK6dmwJZaChLs7vxDottCCqofWq9rSdqHvg1bTpoXel9tUWeWy+W
zs45K+x9IIUu+XbGMK/IxRaenVO/XG0tFgQddl78ntug3zkDXVIPuLNmFR8YbSX9
5zHTS97Gz+T1XjttyDC+wrVhD7qwu6rUFBk3DCKof8oj+0w0ZeRdPUN+w8KdvRnl
+WivqQj3RQwLLILuNJFlpn0iOLMcMZF2sqOzuc3dxc5F2J0yIDgo68k8rthkDHSq
LfnYlE8tRa3scdnRrK5kn3GAp7vIWhOocUSQbA8Dc3jGN0bm2WSh4UYD6/NF2jtT
r/1vn/RXuZCcPPr8PofViyF16Fe+9iPolYdJaNtSfEGVMRbNsCAytnSQG5jMXL6p
7kTu18J0eB5K/5UpePTp4LirVm3OWOz7IvDlyqVVVIfqBM2S7sU1AQH4pkIGHEa4
r8RBUX8xgKOR4WrqLzuhvtKidXsoK+xPaT0s9q3Te56xMgYaZja7KxRFn8TBiH1z
GykaHbsfM5TSICkw1H1NAkDx0O/dBAMGRtR1SKhXVF2tjuUe5Svsve0id5s+zoCk
U+gCc5WJ5Jqb0dplglxqTA5625HOrQ+IRDtZbmpAw2wyE7XD1jq7XoIBeWl//5WQ
HydgEbdNM5jdF4HGTKtH+Y41qQXR53VvjLoIMEp7CBNH9iVhHxWQM+ViIRx0xIPT
sKC6yLZb63YNWTCg3PzSWP7pqzI+lZnSSPgpgE0c0WNBIaR47ZRYjvD7hgPZJ8FU
NHc7uw1+o6pIUyyjYX1cl3mkowEkvqPBtEfD6w4weRu3WhwJYDBsQMXOpL+OtgDd
1SOKmgDV9eI92ojQqzH5KuSXu6IB1lRE+YF1WjuFvq0flV7APE2fS/n0Y6tplSZr
hQhEbmpXqXIfl4tquBWp+W1lAPBi4iW9iYE0GMM2PPp44MHlCdfIxfrwLCN3rTCn
wFZcokOdWvtUgl8oWDEXVhA4T0crcoWOaESwUFEmpr+SjvqV+L2787sG6OmR+u7M
SkcmrXg2khk/0ezfIz5HA9ldY7Yn9GhwPn1l3/ATm17NmIgaqv+IJ31n7SrSZIZ0
uQOlV7V3CIHD8IWbHZVIEN/0pUAwJ5hRPGwcsBxngyyg2qPRL5Pk8OUPyhfT8RwQ
YJ3FS5mP6l8p0I2Dc7vNrtQEozl1ZUcHCsrAjRxbvoWUeZuRX1/txGH95pAtsGZh
Q4NojNRLeUzaA6jYATJTQfcLi3GY0OKi9GWA2i9G5Y8zp8OkOYul30uCEzEztlx3
P7DkjZNVxYL203zugQCY6yncUb71DytUoypGWmU5+IGPL09Sj6rDLwfjz+LIeduc
6oMMtBvUb+Sb9LobHfxlyFmdFM0LVa56MAS6RHV40JaH2Q85ZsyCjtbHpniUQJOO
Ea04j9vDryAlmvuJPhLUxKLkOtbf0gklEXvyeErmoy40SizlSOj+NBR4oxKahqOG
Q/qRJo2mntCxJa4wVkfcJkLRg33ajwDauWUTiKcplYUueUyqpBhFyhuRDsqLCmwi
LPNfhhlhBuXKWXReeNQdXlNl77D+siUIFvFvHBx+VG/ElRSPPbpcYPwjCX1MiBg1
Mvn7dIVpaPsImCFGKyaneHXKFu+cNuW0vkiuF+jNDtli8SjOyMHNSpRo4Ou3ofcL
qpqLBrzCmGqOrl6C18UiGhGIB7tH/KoliXLN3BhqJDdQ9noMn9OWAm3myJgi8SK8
enkfNOaQbN1fddXciR/Znz/ISJ1AfYArFLDZv404GNxKsKySdqkY+F4xc3UYT1YD
PyX6yDQNwDPHe7OxLScmV1uXRpin/IyUe4qMp0QD0/98mHxhVD9LoMNdi7x9GBF6
J53wuwwxqOVOsDBugb1kRwoJZsUrVCDwghpGx/K3VjpK1Z97iOqgx+gOzEp8G8XO
4XGktmGfNl3WWQqoyVwUxwaHO5707iM6OjIzDdFtxulA8moXQd4UyXEul2ADBgUN
yTWCNyLiwNY88xKjpk6sgCreCtMyNRCuEX39AVl8hoCrqEnLw+Jr+sSWPuruseqQ
CKpl51MLoq/G07t3QinPWJaXLffc1s5Hb7cTPwvNVa0WaP8r9tLVbcTmZKPI5oSz
B5BVPqzOMtCr6dndgMSMyMje89unfqcjHg0znXH04a5cy4ctZ7dCnYsJzf3Om/fK
8TCXa/1v1lAY1M/f9lxxnTHTeObfllyjWvXaXTIaYk4743oWSTVPmdy9siINdUaN
8PxPaJtnufK7qJa82X0EW8a/OtObNskn3VmHpujz63/+6fSo+2VTJjaWmNYE+hzu
PRjqdAxJAAouGiNtBNuYJA+9iuajaBMMC4iytRRwuRMFvP5uNtUW8u7mvhgLSbNo
JILlr6LePL9FOXnSFonClUhf/3OZaVfe9zEiczPqz43Llt8rKyA4FIBV45xuE97J
TRAnxWg1S5eUm6vhLAnpIXJl735HR3oq7ieYnNrW3mMKLLxnM6CwEKW1bIIleNQ/
RaOXTPzfr2gMSFGB06Ya8j0pQ5n83RhXNFkF84/iuoSFVR+ypHSLi2NcPpbG7dpT
G33HLvM2rKdW/c2dLdutlG8bH2XpY5p64jhfDHqgQq1tmyFXwvhVa54z3HMbfmAS
7Q0IAlOkA8oEAY4Qm9imXhKcpFbt6E45quH4+xTYOarqXHPbNV+mN3rC6w0mNX+o
fzaGi8lKHiguSxgCMJpeCjFugofsYLerFTkweXn3RCZV2+0vJ2NrpbdzaItkhS46
NZcqBPtAF8SUchvwvbKYgwbpXg5znNAuOMObW8E+A+El01bKLm2pHK+cAwi3910I
1A3ZAtv5q9srLUIzgzi2mj1ShuKc7TJE8OznhdglJg/1KS/xy1/1Efx+w7ElMg9l
0+e/vLgLKbTGoQerPc81MulnkLgvfb6myxBcw/ZBo4UsgkU5aFATFZyqJUe0P9fq
mNwzY+j9F2CRi+u2p+J2u/jd6yt53NKqyF8hTIqr6kwkKTeb//LjgEFfseRPR8uw
UGGZ2EGQunrHO0Y05Ive5QyL/Sped4XEWSIbsQeoJ/mH67Ua4F2BOKobjPN9K35/
DGh7yBsEvDdEr0sGZK1M0Zw9ja0PyqQCxgNHR2utBomlQyqUDuCU4JLeT7zc9v4h
pYDge37zVJPbYDnKTTS49EuulDOrTLCanK+x5iX1CPZ3D97qGlzWdUQIutcWdkIG
Nz+7tedZMO1311oIGBSF/8efqtKPCdh8LiMRS+3SRA1XS/JsItH/4QCW0GsYupW2
ogXliw0eA0y1Y2mRotyDBiF+gsI/FIIXuY0Z63r/S36KmwP2HLLo7TBw1REqLA++
/bwVgvW+3XpGxe2Z98NZx9ABEE0ol/OqOMiBZHp13qmhY79CFid5sPaKrRpAbhph
MVHiNMbLfBBtXZ4c2a0wUBA0kCYQDelQ5+lsMZEmzsbioQUbSEGsqaFAHjYCrA7U
ZhE+Por6xUMURDFWmzZKMw==
`pragma protect end_protected
