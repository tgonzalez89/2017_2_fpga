��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR���[{�T���CK��TC,���:�
&��d!��]9�'D`�"9 S%�aQ�`!�6������V�W�l�a锦E(�\gC�slu�4U5=1�N�m��l�9ў��P���B�@+yg��=�}|֦���ָJC_��IH��9!�"��f�c� ,�iL����^�dB������L��i����l�,9��́�ڎB�|�b�Ș�|e�nĦ�4|/''�~9���o�l)��O/�si,�����S֛�0��8_��%|����P��-Ҷm/�ڈG�]dFn9݅ܢ��6�7B�����㮺�ͯ|��ɹRy���@�D��tօ�����a�{g�sq���`���[��m��/�ڿ6����N��K�K���Q�ͬD��B���������+�=ߖ����#rU6��UN��3H̳�p~�MFڀ����;����d_������Pn�s���s-v���.k�A8���;���me�X�2g�*̊��{����H�䍇���h����x�?��l���5����/5!O	$�����`�k���4�x�����Ĺ߾�r�"jF�B���w��3V#�􍽦�e�^`*�=�XJN��N��h	B5���B�N4����Y��T*��Z��c�1�:�]�+kKu/l�c���}�N��~��� 3���f���)�� ^��o(�^N,+�V�B��T^NY�����ô���a���{����F��E����2�,U.C�J�KJU�b��P�%\����J�qb�.y% ��R	3�^����(�){�~�C�e�AHx$�8?8���-7��
]�~��`�6��Y?C���ߥV��%�#0L�}D0��J�"��K�cN���B�{SC@�w�}�ێ�=��G^���3��w&���9IKI|5����P�TD�cI[�2]�1~�/����P]���|�����z0b���j���(H�J�H��(G�o�[�´j9U|�mg��'~��-/E��q��՝�*}{�}\ �S�Z�E�������Mǌ�A0�;�Z�,���s`�=c���UV�ST�Ù�+�?$+b���CPQ��G�tc��k��A���c���2�A��j�)���a �	�����u�.�<.���:���1�D�e"������/5�W -s�����\�h��gn��_��c�(\D[_5�8���3���fi+fg��S�C�Nl���͂S�Î~|S����Zᐹ����4;��R��Q=�0{ĜG�����1��,��Թm �k`�Jm##OG�4>������@�M��w�@��i�s)��#b�]�&X�-�������_��|N�M~�R?>j���b]pv@j�I�}�+�=�`�{/�K�vX=^Lg�<�.r8^*��7���i�I�j�X�n�g� ��C_N`=`��-$2��U ��_^�1��#֓�8��0�����t"�V�su�R�u����s��b=��ꏆ��G��F~���G��Lh�<��+����z��XQ��1�-�w8��I�j~m7��2x�'�?�Ҟ��Ej����m�TVs��� 
M�.���`حqk�wC�f��Ά�O�K�F��|��bj���O��=�,/CX����������-����t�x�r+�`����������.� �Jv�
O]��׻��L���> �6�������l}���_���R��8&����I,�����ኺ�{sR�^{�����M�?b�4fq�f���e����BХh$Q�I1��*� �ފ*,�oH��1�4�/QƖ=�YY�.�I�KF��
��X��Qٲ�X��	�)1N�j���om(��ꐱ���$tm.��.����L�_�-�����-ebn_ssN�fQ�z>@R�Z��(�j~a�	�1�.mL�F��>�g�l��6F�~���L��bYc�vY�[�<+��}m�I���7=��a�8��8�c�U��~Є^t�ݰ��m�B�n��'Oȓ_YL�=hGғ!�Z��"^�N�ې?VI�Z���P�Jjrz����zr���I�u��d�ק��1FX�FO���K~��B�&��(��g��;S�=�Z&tM�M��c�@�p�ć2���r�ƿ#������iI�*�,����B�Br��C��eӳ��H���-B��5a8�:4n��P^<�
B�����B�~5)�C!��8�J�<��H�\C(�˶a�K��v?Ҍ�Y/�����g@�u}�.k�7�o�;C.�}Ζ��uh��Sq���{����:s�m ��Y�j��A�']��'�뷱�U!t�oV���N�P"�����Z=+Y��c`�b h	����Lt��Y1;-DWz�)nq�o�~���A��E�L7���4�>�+��}��A��h{z�/򔉛t�fgJ�LB�c���W���IZ���\�S�Ī�����tM���
�N���,ںuuYl2���b�#���I�;��!���>!F���F����Ø�W<��<�9� �n����%̭��?��uS.�ut2�u�_�|�2�7�(���1���c�o�dz�p!���c]���������Hn�}W�`~�҃tF�W㲤��Z>�֟VN���6�S)d_�0�����o^v����K)@���~S3pdgv�*�c�+^ݲR/��J�¼ނn��(�w
T"�/�7���F�a�V~$������J�+�ĒivdϿ� ��38�����m�N{�wo`�>0)���DٜDI�ܤ�5��t���*
H�>T?�}�Yye=:�U}D��X���q�&D#��h�G'�z7$����g�e��e�a����\��l9ȭ�����A,d�r�	�2~`>r2M9�eL���l���N�s1���w !zP��VV0 rE�Y��Qc�FŜ:%�)�@��#�poE�����s?g#��ql�O"���T#U)�>����ٝ	�"�%���˳˽̺u���+-b�Ԍ��ɢ�;�-��,	�i�,��0��E��n��L^�a��]�g�^F~H��,������;�F0*�V.�r�{�y��(�eC��E{�f�AvHm�����pn�����Ζ�G�3$XT��J�����D4Y��+�;E�e� KV����Y�ȏ��L�����	�*�G�AY|����X�w�7���X?�%Ԯ��D����{�E�m��톘�V^��gŐ��f��sa�b8y���h�h��n�핋F�E�# ���ga����a�@NP��m�������-���03���׋l�㫢�M@���Oo1��W�F� 9~d+;�P)����AO�����S��0�~��_����MŬ� 3��Q$�����m��8����5 ������D��6��){R��eݕ�?D�b�}^���a�� ~���bE,{�Җ�������&	Ր�F!�h�6�;QY�@R��Y�UDW��שrSE�!囔�?��oZ�����3��0��v������0x�8<���3[{�TE��� �������u;��)AO�Q�mm�<;E�&�G�7�������Ú��;��r} �����T���i�΅���3C҂P���_�<�8�D�N��a�!�ٕ$X�{ޣ፰P^�+�x�.m,�%6��nk�%�Ȥ5ɖj\~�\�a�Y2aL�)K��3��B�+�?q���*���툨��~�J��5>%ÒYwӑf������1�� ��ȗf[�H#�)��eW�/X�pQɑ�Z׻򈅇H���5�n*��V/�{LJ��A��L��C�\��#Fr�H��ќ���2�ˌ�Q�~�Hi��G¯��� d��m�� �g��"��$d����֏%O��1Ӑ`�ZW��9[w��k�[Զ��7��%��ʼ����*��Q��W>���E���v�=�P�}�`߰5X���2t^r�4F|�(~�>U@Q<B��h�4uj�Cx���q$xi��S�*�S��F���O�>�,-S�
�m>ɹ@���#�f�M>��ƕ�|u������VK��]���KsR�,!�o�Ņ	�[`[v�"Ȁ�`��w9���0������m��w�W�h~l��)���~���K�tJ��w����7c����Qɬ@�g@֝)�n������YK���������#��^��Y��@�md�p+ӈ�s��n����ԜfG=�����5��U�A�RYg`Κ[���g�� է\��i1h*"lsm\��}���9��RK���<�:<M�[��b��֋�U-#������"��	O=#�g���q���RS�9^����ϛ$��,5�QG�/��#�)"X_��6�k�������z�:��ݔ�̠gX���zM{a3VˣW2�H�8춞K1Z�%�<8e�&���V�L?���c����tz�
���JN������D��5�j�Q�5:q��( ��<&;�v�f��B(<��\ ���z��&:�����Tm6NN���wì������+ g��j��vq�����g�TV܄�	��73�@������-jീm�d�<�]�/@Llј�2����JTd�`w���ƨp�U5]�g�5+Z$r��qcpoq�}�
�/J+t��E�$sEpE_�:���o�'���^	�!�nlF�W��k ��j��K��	=���n��l�|��G6�}~n�\���7����T�4ـa��x�T"_��a��� Ef�W&��� 8�XQ)�K�L�Hܶ�CT�j����n^�o�R�(ڕT	�!�jDsN�O g�6~t@Ѳ��A�1�j����T���BN!��fJ8��/���<.#�Ͳ�I^�7P1eg.��}���^����0�S��ta�r�l	 :���~M���Nu6��f'Np��9�N �$�t�r�_�p�������_�V<� 6�C�9SF�*�]4��m[T,�D�����1�:s�L�UC��~�z~Ƈ�0�jd�b��r�݇���]��Y(���m��g� �l�U����j�5D�i"\�ֿ�l�O��6|�m4�hoI��b���6U#��&�\��v� ���z�����+ǐ����AL�(�C	�ךQ���i�����vu���Z;_2}p����	v�1�^̀^1h:���� ���m�Ed�+ڃ\9�!�H/���)X�T���T(
��jRPC*.X�g����2��\brW~�(�i�\z&����M�ه�b����͆�T����RF֕�k���]}r�nٷ�?.��!��1�ʾB$0y�u�e����檤��'��!���e�1�)��p��?�FX�U����>n�%1�}u=��+*�׽��x���$�P��YW��=.�"yE���? �̊� O�lo�$����ý�^w߾"~����Ǒ��/���/�b����^2�-O�44 ������Һ9Q�7N�R_J�xUW������|gW�_�ϥ�-I��=,[�'�'fx4�ޢ�R+M���0_��Tz�!��?$]r�c��O�����{���'G�Gሽ�1G�i����s���nv��Z]���7�k�ވ�9��+.r!h���!���Ӿ`����(�+h k�@ĩ��[w����w���v��L0���{��0}R�+}��_��S+�~��e�ϗ�3�M��Ƨ?��dr	���D�s�S�)���K���q!B �|���<49��͖a}V�=�M��4Lx�5S���s�n̅�Y��M/����7C�v''����)R>SJn�w��l�q��pؓR���/������;5F�@���QM���}^3�-h�nK��]:�+��2��� 1�₵L�J$�� �˒UJ��b�a��n�K�����n���0��D�h��p_͡�}a(�HޤT<��G}u�k��G�������?�爖}�`n���YD�F����;�o������to�Ә-^ۣ��J�ͻA���V\n��F5��7d�̳8FJ�a��r��$�ʁ�He�r�IF�s�K�B|3���,;v�u�2cq����I�Fo�����%�U���v�|K��5�����R����ͬ��MQ����!�}�]�?�Bڲ����N3������p��;��<�u�`QI}�u����e�[#m,�Q���$��΅V>Cm�Dk����~�V�@!���р�ޙ��&��
e�I���I<pj��&SYD�uB��f����
$�)6!�3ĩx-;��.�v¤��Pd�A8�l/L�c{!9Ơ!��7����8b�SI�.�P�h����Yg ���X��F[b0�)�7�^�4�S��ՔCW�=�nu[ۜ�w\�TY>G���`-��.����>�P�a~�h&����[����x�������V��{e�V�g+�:b��Dx�=\Q�z��lI��l.6V������@����:Y��b�g��@�-�����X~F!������\�0{֜U3&��;-���21?�{0t�)�R?�hO��*Ktdi^�fD���u_��*�R�d��{H�l��yl���!��_�pyS	�=�b���~�F,ŀBG���!WIZ��2!��X��4p%*E"
��r�������a��*@R����\O���
���C.~�p��
%��{O�9��ե��Ƶ=�
L��c� /�ג���_q�H�������e0�kmf\'��<J>�'(ϯ����H����!�zJ(+���<���ʩ����b�q��L8��pΚ� ��z&Z9�(皘≒��Dݎ�3��x�L�8�_a��y(q%��wS��0X'!r�<WQ\����H,���}���������7�����h k�ꅰ�����_�<�	���)~�k9�/7t�e���9�GK�@G���t7v��M����l�;�:4���>�1���dNS��?��w�x�K��kЮi@d/�c;�8�;�A�&�{���w0X�q7��Q��H�ybyۇ+�Η e�ga�#�F��0�Ni]��]aw8�G5��x�=���뤦J����R��rI�V'�1V86���o[��~�$��ևb��w>)���{k�`�keͷV>v1��j��:�)6Q���[�L�O.�ߣ��.i�o�ڸ�X%pv�L����r����Ϻ���c�	�3W#D�EϜ:�s��I9Cn������}�r����F�1-��� O��LD���2�7�/����\�~m��[�6����%M3��
뫝�� �����ƅŠ0t6�y�O�x3� ��N]g2x��p�� wLAb��]>	��	ӡ4\�9)(�t��|\%{¬"��F��*�?�@�M��]�	>Y/�/�|�ZtيƟZh�{`�leˏmC������N�A�	�v[����m�'I�E�)�Q2YY�LjUœe�쿷��K��j�&9�!n��Hiw��Mj��7��4�X`�xwb��_�.xn�b>����xx������u${i��˿E_�OR7D5w�*"hG�^�8[\�{��C'�%�6k0Yމ0�����3�LC6�(��vm�y�3��Z�|N�o:/lޭ���'wN�����-	�LV]@Y��R8`��`K���.P>�(�<�Mwz�cD�U�Z���n�~&�$�j��u�B�������a٧!��	��%����������kp��;��v|������ǉ�U[���ս���C�&���3`�(��+P��e2�&f��sW��σ�h��_R�Ng�2($�Y&��}�A���6�����?՜\p��:\�&�I)���ĎO���O�*c%i�,�\YW��4�#�����p']9'���J	hm��ݭ|���QO��֢P�9ȸ��=�͌Ѿ=��x)�ѹ���G��a�0[@(G-��/K�)�>&��Z)�ߟW@�������[[;\]Hh!3�B� T�}����`c{������cW�.ܮ����uds>S���.���^@v���g$��K��Yk���m#5X�,�^Vν��x�9+��� k���q�"�XfjW��D���:�x=�S�Pvq��Hh]~���0���N���ӵ�5f5��2�#ު��A-�6:&R4.-��@YR�?�E]�~]���;|�E�Z�^\TT����hH�Y��
c�¸G9F�۠��)���n�R�[窷���Q���B%f��J�8���|b3K`���O��w�I�HM�/s�����r��ydwQJ��ją�b�xwLۡa\S�:wWzPQԞ�Q�k"������p�3A�es�?Y�n�e���;�.�ؒU3��#�LZ��>���
5���5�I]&���Ů�	6���_�⟮�B����=4�������y0�	^��@i���h�/�IZ��JW�`@Է�x�ϧIv�����}6g;�?�y���ae9#�Յ93�x|�tP�S��+�T���g@d�yq*y�[��(6v�K|D��,pȸQ�L�Yu:%{��R���-��z���
���M��N�"�q�f��ez|y�P_g�]�[�φM��ł� fR��=�Η>f��� tڞ��(�4�U70�2	&���u�)Rb��ʯN`�s�����0�,�0T�  :�����{�i�����
�S���y�[J����2
����&D��]��r�(/mK��^-��.�n�)ku%^��H��zݨ,��H"���qa�Q�vo+�y�Q�Y�x�]13�?�Ar��?��e�D$
t���L�Q��˃�OM5"�n������p���y�hmYP�/2�^9SF�B���i8�(	� �~d	}2.j��>�@�мh�񎡡8�ׄ�d��#������ڛNg]چ�k�Ͱ������:���q����+i�蛠��H5���A�G,\�H��*-Q��İ�j�6��nI�b$}�&�Wk����,����E�=0�']txFgC��VM�'��j��/9$A�ʽ����Y\�
�U8(2ك���T7���8`m&@>3�vH�6|��v&���C:wv0]#����_}D��!�J-�BW�M���ΰ�Ig1�;A�@!־���V���w�(7��yۼ(�fâ̗gM4�Q�c����$v��_�"Z@�V
�3e�5����B�	?GF�#�ǔ�ۭ����b/�dF�5���~�$]b�U?p���گb\�����(����Jj2�cP����$t��b�C(��R��F񾯫��Ԅ�LmXP��$�`��/�����怚�O�Fm���&%����+?Y�f3��d㭜9rs�Cg��Z���܊jZ�>s��L>���QZ������#\��w'�rr�����7��������ң&�#����=��R���H����PU����v:ZQ]�lX�@��YhQ��1��;����00щΠ�@�DPI�0��f�~�,{f,��o�R�7����,��@u�t|+ToC�}���,�o��39�`DRT�Gދ�>�FC/�6{�h��:�6�R��$ۖ�����E�W��1�IR� j%U]K���D�NV�*Iگ+TL�$m��fS;�y漂�;I����UE��A�k���]/��U E���U�*#�/��`��7���:�{j��T�E��w�������o�YF>��&׺%����Ӵy#M���d
������j�o���������!�H5��ҷ	wg����T?��2��+�M3#8���_�^W����y �ΓrX�Q���Z���ە�f����R'{��'0h_v"��K�I|I�h�H��G6X?���0$3®8o2�B-dvC�5;���&��_BM�9�`\�d��o2Sg�B8p����������D�6�L�ڍ7�:�q!�ń|F�.��� �SFݸ.�KR� k�����lm/���}B��aV�l���^��a,�h*PQ�|�V��%���Ph�\,g_	ߙ�q�CD.z_��m�uHx���R��5�ĦՖ��m��	Wmp�q~�_s0+���SqP'S��g�Һ�>���D�����B��=A��3��ǘ^����گ��4Xi�k���ҸS׾>�,��0����3��0�q�����j��f�^��5*d��f���\�6b�	&7�hk)��]��7|�J���$A�I�QJC"g��Jnb���˄s��Ս�Q�n�i%��m�cEQ">�%���ݏ/t���3nG)��PJ�R�4y�5��T��$���,V<v-��)xl	kLҚ�t���0�v�sH���		rZ�e�~���
7O[8k�Bg��CD�cL���.Ǚ��b�aR*.��T�Y�;�ȍɄ���Kt��H?�k#_��ո�Q�{=z�Vy�rP@չӌ�m�G �.����!&���4��9�'�H��d'�%k5G��71a���R-E�?6�Ľ'l��l�a=Z����s�D#�:�#d�k���c�<x0��pGƳ�nn:j��&.
�'g��,�W&CC�"���/��K3��6�ɄS�h|k�q�W݂��o��Q��H�бԁ��D�K��H��ǂ%��jm�� tUK��=|.Q_�����w� �	�7�m�o��t��a��t��K��q�bNdPnA"Pj%�~v>z!M��xA֧Q�ҧ�44�sS��z���r��E��"g:cL)��<T}�b#�l���M�+� ���U�U� ߔ�TeYם�/]J�ޟ��Ӎ�ɶ��A���'��]��<�Ӧ���a8H�V4�m1M�K��	l��H�J\�ͽ�#g0���4Ҕ�J)��̆!!�,�S3C�J;���B/�]���D5����v��pEu�g�=�&�z�"�ۚ���7�=}����
S��X[�v4��݁�C�4�du�)�v�uC�2B�����M�0�<y%�=<2�k�F��"r)����hO��q�t=�(���zs�2WոYϒ��蓣��vN��-���aHM����:	�5U^�o�S
�$5�9<ҰB����uW��� �?ۓ�K�>��U�km߻Y��&�2`��9.���<�p�w�h�D�,��E�ĸ�_������U�����-�Y�����(����4Bا�k�>�+�u��¤�U�)I(���j��N$�d�]��E�0��vn�Q��K&��%�6o-w7�P �E��	\α6��P�5�QQ%����(C���3�����3���C���C��v=��:'](�h��ǤFJ,|�"'ۆ^X�	���_�Ln�$�<lo���UJ��+��7sP�����	�ju���}r2��C�����Jj	�����T��U��T��~ʝ�G��y!R�Ko�`8�"��t*����pcS�K�� @2�s�A�{ͳd�������,`�e������{��1��P�?�t��p����H3S2W�c��A�|m�9B�U���;�Z��ȝOvV6}V�U��+�ж՝��<I������+�>6g��#�.�Z�˶��/t���)T��΋��'�9��=�j��L�o���#�����R��$^:�:�V� P���������̜:����^��G/9�(~�Q��uy��<F����ш��l�T��i�BJ����])^v'Щ��SEi�'~����yEr�~��F����>|��]\��jNɻ�Ki�N�`����V)&\���s ��N�f��?h�~�*^g��޸�ѓ��b5Lb*�^8������_�mW���tx����� 
6X�:��7Ѳ��2�aib�
�iZ.��r9ܨ��ʉ~{C�bC�b7Lh��[��>�2�PN����n:�듽�W���o�ݾV>J`�Ӷ�#���ͻ��#�_,�weq��.ԣZa����	C��ך�My��" �_F���A��	�^��<����!3tQ����#�[�>��SI��b�	����fI�c�i�m�<e�u��6R���KC�PdɅ`_Ջ)O#Yĝ>�س��[YYr���γ�A"�'����E�pF�t�G�~�1na��/h�h���	��H���#�i��v�������	������3��r�fW�vej��,WV�ly�F[NE\fe��sp�S�ջg0��C������x�w�h��?�û9�_��V�l�8�r[��~��mI��]0sCˤv����#U��NL�N��`@���(ã�,�ȁ�ow����8wp�u^����^y�9̇��ò�wC㺾y���q?ve��� �ng4z�����V$�d84�;�MBx�g�a�N`&��1"֫ӆQU�G0�ذ-���al3qrm����y����TxU�㨈P��:3�Uޟ��D���#̘_�Z��}к�1�a��&��Z�:���<��MM�\8�V�F��U�/"?/�M������a�x�*x��k�K�S2�n&+PV�!�������w��x�b]?%��(�ux�!0��S���4�)Z��)�L�I�o��7�u��:�ʠ�XP�z�$�g�9G�+c��ЍW�s)n�0��q^�ú8b��b��1z)�)|V��s����k����!��;�Pc�eI�	4o��58dɪ�{ms�F��87��&��7�<+UFD�����?�z+��⥙�p�B���@�v?�K�}���������
�z��Q��������J6);��%j��ſ��Fj�)X�]u8�1F��q˳�ȅm��(�2ߪ((�\�𨁛�1-to�����/���A|���)���%�g�ij�h&=45�\UC�l6��x�<�vo�����!��8ʙ>�č�r v-_lwIlޖ�e�B��m���l�Η@����\��80�u��_�G�'��kI5�.F��� )M."C�Y}��j�=��-%C��W��k���qE� �z՝8LO��'2�q@��j����u���Ww��X���щ��!J	��lHo�a�ۇ�|�f@�+}Ća߸�^]6����"�>�^H�R�3���Q#Fˉ~#.Ds��ԔBwWK>{���r�4*վaW��	��{g��1�	����
sQ�k���������9�{�t��1Q�s��%۝�;&\)������G�6����Cvc���W&�u�f��GFI��Cp_y��Bef����8ll��(�P��y�=�=E�����6I�"�qL��i���Ï_1��OsS(Հ�L&9�fQ��%�¨�OJ�f7c�V9��@���G�eL��K߆sg�V|�i�����~;��f'�ſ�݅f��Se>���^�mo�0{��馲�?���pSWH�ٳI�UE�!8ƺ2����� ���*���1u���F�p�Q��W�[��S=�'ם�W��'�]�����c���	aU�7�O��Kw�)���5���=�,��>H�$�Su��x�1g+Gm?_���O���������^�p���	OD�*G�n~;�N������#��a�8�سs	��5MG/�8��k��M�E�~��U��|��M,�O�
n00�n��O||�� :�8����J�k�`�)�['�'t�#X֜r��������K=~���Avԙ��*���%�be[a�Η�4x��Q��z��F� +{��DCa
e��j��e�O����R���p���P�N������\jG���nW� �O�;Է�8�t�����f�;{���k�+LJ!���SJ>�Pj��gf{�̑ŉF�N91&!��s���ʻ��ǝ���� ���k�7�9s�������@b��4����Q�$��6"ov��,�P]kqI��q7Z��W)�ï���y�����P�R >C����}�ܰ�f<�3�y��a��g;p���)I�80v�I�5������ӝ��a%�����"��v{X��WaR�U:B�G���������A�n�V��vu���QhBf��:�����S�M �Y�>
zj'�?K߾Y�-��� S��=����r�~oM�����z����PĞ�(�kְ� W�]L}<��q��^�"��_�	������3�����K,E��n'��j3��P���ϭvu���&�'!�0ː�@�\���*��+V���~�Ɏ$��)ys��|�� ��"�!��
��^���:� X�8w*qwAm%�G����Ѣ�B4 ��#s]���*�,�C(~�%!��\�D����;�WȍV�ǇϮ.������\���q!)��Li�
�5V��ԡ��dy�>�:�8��q�rυ9Б��V3䆈?���c<�~t�o���	G��ygn��v�.W��@��M�̃P��9��T���	�������άtN,S��K��b=���gZ��
����25'Ir���%�����mC@l�m{�����	�e�dRR�'4�M6s��}�@V�*D_���o���g�9�a�9y�x��艡ݓ�hh�˩k6>Ո��!�bՐ>X�+���:�	d!�"/�ݡ�<#X���Q�zx�J��׷;�`r�\iuK��9G�9H���Jb'�dQ�:LCx����Tt�Itu�G�3w��~��G6��&l���������֞��4�A�����!��/;%��!Nzf�jE��]fs1�|2�D-��c?���~AS��Y�@���]@�*�U�èco�͐�e�;�{>1�<�͙C6�Qo#�o����Łd��Jb��W�d
���ݏw�6�O��^^�z	�#����@b�|Nz�#Q�k�6YUg��GE^�4��>5a�s{�$L��N��$۪��7
�(<I������� �G�-����ǅ7�@�К6�j�_"|�8C�џ��w�썷o��S�D ��.�H-PA��v�3���/C��E*-�d�J��8�����Fh�op<�R]���?���i�1�A�Z�'���*��M<�tc<}eZl �µyN;���<p~��߄+W5v_�쨵�F�Cmz�q��J�%{�F�W�N�EL	=��td�3r̗Ta�C�e����L Ms~'���(�=�y=C�_��*�S��F{�$`kn$H���4�b�R�� �r��t�?�&��/�1��a�QH�B_��u�Wp+ZՏyŵ8I�[�a��h�2@�Z岙�3(W�C��~�j�n�Fҧ6^n
�߃�)����C����*0Ks�e�$�G%��t���(&}�]n�F7��m kn���NR�������ܟ++�Lsx�z����V�E�n��H4�����Q�>�7��ޢ�+cb��=(e�$��'�Y�k��\s���ȟ�$T�j�^w�U8� �$��waٚ���U��E���%�@N�>�[��wR�BW��i���(�@B��L� O�������%{3�Z�S�D���]FgVx�Hd,9uS�ַG�Cʹj��;E��(۠�ƛ��)��g���0
\��A���*�Gی��Y~:�1��_W@Fk:�r���no�3�!���~>V��H���`Mц�42��W_6U��iwiig�����k'�E	i[�(Q�,k��ޡECx_��R�-9%��ە*��
9�w��~�0����:�@|��NG��;�/�q�"�h�崃�C=e3���O�L�~����� �ܝ�7�H·@� J�OZ,�����+�a��}�X� �]U-��0�狀��!� ��hw����t�qQG
ݎ�fE�/ҏE�q�h��T�E���j�%��BA�s�iH%ϕ���k�C���2��2�%C��uVb!Q�N9�^<=�;��h�Eb��������&'nV%uVT�/��OV��������L�c�c,���f��#2ǝGa"�QΙ+�͔���kT��als�*�@�L��50o���90U�ڂ����]���6��W�:����#�I,�w^�-`��me6j�ٗ^{�_�{Jʓ~�t>MovBТ�,�;SՓ�F�Ӆ"�	?H`�`b�vQ6��tgT���a��E���9�.Ar}:8�����-ِe1�^���wq%˲�#� �ފrD��舂��歷w�t���f^���Ђ����p4���\b��'-�ſ3�`M"�5�Q����NȟZ8�^���Z��t^���>С�HVu�*�����w�}�r0�PX-��B߭��֔0�߯���*�����(	/@�طC#��������m#��U'�K��T���2��2T[��]o~�פ!<xD
��8S��|͞2�Ө⶜�T_�+��I�2yJ(0�̇�B #a^��S7��q��cSq��̀������Pw�$%X��ݥJ���3	�Yd"�`��j?*?��j�+V}�8rU|py�����%}T_&�0�����<��7��	[���Ռ��H��1��0ӷ�V?�ݞ
�:!L��,��2�pK�Ǝ�6q)Ӭ��țF�t��\��u떎Δ޽��[4>�w/$5��Qr*�Sc��y�^c,Jpu�-�d �M8��K6wֳ�ꊷt�/$�S���Џ�(l�>A��e�ĢE�����5I��W�)�˛U]��![�Mw�x��`Š�U*��=x��VN��0���<�	�x�^5������H�rj�V٧~���y�ĝRӂ�O��տ��c��\�����e~����P�Ml�f�� �gD��T}�G�Q�������̴T��ү|b����g��!nH������<s�<͟�{@�hF��>�Q�+�;o��f��l��~�Pe�	����+�~C��)U��a�	�B'���ɬN�5�V���ܫ�G��$ � y1Y^�yB����ָ(3���R	;� =>�:S�3i�L�_�z��#�^����u��:�PtU/��[�.pD���R`��,�|�ݮpm��8���y��/V:_�Uil�Hؿ�f��Yrrp�E��iX3���Gc|�~�o��X!���A���lO)�2�n�։�׍D�q٭E9筞=	�n���{�Qӕx��GA��0d��K|?���<�="���ǐ	v�LO	��e��&K��M(�����3�j�3'��s���ϕUo�X�G��ؗ;ױ'Û��"(����HAǁ��㇫����#v�Nɯ�j���a'��|��$]~�D�lH'��D� b� ���D�%�Yk���T#6'�����L�0������A�G��!;`t����9%*+�{�7?ge�T#�r�i�ƃ���+����y�:���	�;)h���G*�ο�z)��!�[���?iY�:ߜ�~�;?(���e�z�-(�i@n?>u�Ľ�;=�G����vBIgk�5�������X�O���	�����	, cT�= �@�#�h�9�G���,OP绤�B�*`}��� �}�m((I���)k�,�	s��7>�3B�.g���W�y�����B�@�2�<	T�v��l0G�ǡ+���ٚ����."�q��(u�I��ZVo���Sk��A� �F�&?�Զɕ��S�]I��(�����j�˿�B� oP�*���"����#��=<��nД������W�6=c�'�V�߶#U��rl�Uʦ�:[z�{M�Ҫ@v�i�\%�-Js��:c5fR�V�R���#������<.olz��ꁒ��Q\<
!���Bߥ2��4�o����Z�`����h`��3�(�F;�]O4n��!.�r�ae�`�M�^7��ȉ�aU�w�CN�	�(��N��ms���<X�R�2���3/ږ�����%�����K���:	�V)9�F(q�j�H����6?��M��zZ@M<��`�y\|�ڃ�3%�6]����9�o9���;�(*ku3���jW{�՜����{�H*G&�K��`����f��i��}n���JOi���@���ҒJ=۔-݉��V����0���$�=
������o���l62���W����-���l������/�;3�ޛ� ��5�GL	�
)����.�.�����3���\Ѿ �|.�ja���̩z�/NϨ�����]1��0��j��D��/��h�{�����i�������k_.�"O�?� KJzQp-t����o�.��_]7�~�FJ�M��B�S�a3�B�h�T�
/�!J�GX��+��-h���.����&9ٿj;/�����������k��a/�"t�?���ՠT�c7�w��X�ؙ]]T�ʣ�0;�7�da��gw+����ς��C��0m��<h��zX/���R�TvK���:��W%���1�c���N�M���-8�� N����ăǯ��a��pLk���n�'�;LB�f������T��є�n
����XJ��k��������O��8Y�=ؿ�"Q'�g2�� FY0��=IᏘ�ƻ��Ȓ�-L�Hu>ӣ��J�]�!~��jqz7���[�kL���]\w��.!p|O�Rqʣ,*�t=�s���I��v��@/ J�o�,����j�%`�״vX�f��'f�P<����v�&O.'7�U;uҰ�@`�p@R�&��2\r@!���8`�M�.]��jf�m P�Ɔ7�W�C):�f/[�0=u¤s�*�T��L�l�,�� /-|���/�q7uGl����yiEsW������<����{aSL�����$�YPe��TMl��Gޚ������iN�k�[���H{6��(�`�Ä�1�+YNu$���z����b�Gv�K��q����
�x'rDLY�P�"�:L�$�_�~��$�4��t�(�qƚ���s�P7Io�V��iJG]��zƱ^�h�����m�8ct��n�i%P�l�ٴG�"
�c�xw����)��*�����I3� ��[�e��+G`�O�C����N�#��?�~[��)�~f�x�0~�z��v����+իr�d���y	P���nn?5$�9����d��s��	jM��:[5Y(�&f=�%�eM�v��{������$���M�Ld^�~"�
T��N�ا�Zu���D
R��`J�$Z4�6Om$�|�����&;��G�P��W3�8�{���b�������_����ňʣT a�a�Zv����^_S��L\C����<71���}|�u|��D�\]em!p���}#[Z|���:��Wc��3��Pf��%i#�gL��'��-8�x�U�	�y[�,@_A6L�.���S������Jxn�n���ŵN�V2����қ�)W�lK��"9�E	��[\}�X�c�JS�T��p޻�4���`��u-1ρ@�]���?�9e�*Z�$�3 �ܥ�5�޸�R���
)��qc���n!���V;�W���ǫ�P����c.��K"��@�޺��$�5�P84v~GX��C�NAl(�V�u�$'DBP���pY���2_<�]Y�!��H�l�9�#��]x	���`��>Z��	�9�b��X���{�/*�G�MlJdO�Y�U��4��p��`����O�lNB���"���l`���WDY���(����g&����>%z�i�JP��i�D%����b�����j%�Cg�#��9�j�����x�ۀ�u�[:,�"�(@P����:�4��@��� �ڝ�}��x���#�S�^��%c�)U� ��	��qJ��B5W�+�K����Dh\�v8��п�������xW�S��2]����C��g��:����W�ڬ��M���	w��M����H�-�uڍ|�%�Q��<
N��1�>�
��7q���PΡ��Sjz:�\Q������G���e|{��u�7�$W�L��`%G��y�i�1�q�7Ρ��;�X{R۷�k��Q�LL�����~4ke����И���b=�nm���i��5Y�gI��5�fv�_�*�@x)M�w�j�n����H�4��N[}�}|���_�u�ğ�y:;6����<7�=�8�^I�(ī�|5��+�h��ɪ]
L�pՈ�����V��t-E��*�I�����p
�e�^��K���3	n��=F}��Ց+�ᮽ����s4λ{�=��RI�ؚ'O���e ���������<�S;��THhZre��bu�J�tͤ�,�^��lS�l��� w����m���<�؆.}����k�UֿH��CZ��v�{:d�k'����)`x{�k옔�dy���ܛDRY�O#=id�#r����.�I
W����0����2�E��(OB�*��qte�q��|��al�8'��R��2��SA){�n�2j�Z%�Dy����-޲�W����� �qc����J��+��vO(�b��r}�4�/�1H��s�k(��3^�����ϑ^5�G������0^~�ρ���m*N  ��.$�n:ө��5�,,q PB�Y��+�G���X��B�� �L�gb"�'$�	��,9j�l@G��9;^�����v�ՃșS��횭��i��g��QZEdټ{�������MX���m�|�j�X�T�O�)!�$����?����!Vj�WlBa/�0!���e�ыR�r�r�IF��s�F@��Y�)'cT��Y�Bk�I���x�K}�� BAi
�=S�������U��]�	Չ4ԣ�|$HB�3�&L�qi˞C�)�*V=�"�֑�m�-EMxȻ��=5i�����Ȥ�>�'�H-^�0F1,�;%J�DE���F�4	��,�)�DQ��{�8o�5e2>�'�,��c��,�Z�*�-��q���ПE����TDm�˴z���i'J�z��o7���_w�֖�����Ҵ
PXuSE��?��]�Ԍ��Yι�-jˮ٧��c���b~ߜ��1�l�*����ZŬʌ���F!���Z�� �0����»k���Ƙ�q���$���0N�'�f��ֳ�������|I�dq��ކ/I5B[�a,V��T@�$�Ȭ�J�������!� �VA\Ջ���K{�"�҉ą�X�f��f��r�*Z��4�@C��Ə������@���i|X��D k�i�@]���	�����F.#}��kA�Yj���*)5}0�^G��G?�+��<����̭4A�KL���}��S������k�u�6��ʤ��(;�d��?��V��O�g�:��Ȇ�[�v�=�H+R��dD�aj�wP�w0jZ>�v�	�|�.�+6��\�@4��,�)��GB)�#�Ae��ٰ�W ��~>x@��ࣱ5�f0�[��m�������:T�Nrʪ_�����h>��b��c	U��ߨ��A$���_|��/V���H��,���K`�y"4��|���0�"c �^̲Ԡ�8b��Ϗ����8
�+p N�}�Z#-�m��\��c8�����A1ֲ���Al�Ww�����D����
-���-Wc�fg�~�����c[Y �Y	Ӥ���&��4�:gw���i�ir��޿�O�p�Z�o���>h�6M/}����?��ެ�j�[�y�W'���"���0Ƭ6�N1bN��4��Az�bݐ�S_5?n���g%*S��Zrw��~A��t�G,Q�Š��{ܸ�1	
:�өH��/��hu1P�G�h,������SC�w��r�h�F��($�3��h��s���s?��\%�b#�tY����aD�p��5e��4X��%�D@&�)���t���.7��f���04}>F.)��>��9���
��%�(�<��:�F���K�T�L�������뎵�O��3� *ŗb��>*����a�oP�Ӵ�+��	�n��{�"��:N\@!�V��:���9oǷ��Љ�a�nYv�Q��	*�����b+�B�4/YŃ�{7��{����<JϚhZ��6V��GjU�#]+oNnc�$�3��.�Ь|�:B���w@�Rr��E�6��-��{�,�d�r�e\5ۃlz?���pމ��x�B��~_�yE(�K�З�nt���K��b�rU"NE6]p���d�$)�����Hℭկ;��>�J�R#� �#[�{^<�L��]3̴^hA�г6�e籣Ɖ��l���o��[(d��47'	Ѥ�.����ifAᥭP5fAj��>�)�5��Z��]��'�&\�~�Q��I����T�T�i�6҂���ug��E�^	�̔x0c�_�Oc��2u���HA'�B���B⽉��p��fş�6Sz���=��r΃SŰ�߬���ܨ[@��-r�Ǎ>�pY��.O���~=)$���m�Y:��������nE}�)�!��O�S- Hd@|W�.��tTu2 ���Gx�?�u�f3*̊�ۯ�u�'(��QѡGy9+ͦ ��X#�4��GJ�@V����uY.�T��K@�Q��T1#	f�Yb.�t�Q�:yK[�b�贈8�렂̵��h�dd��HY�ǻ�[�氙��H��&0���3I"�d���@|~qA8�����'`�בJ��� �������ՙ����W�����~t(�]��A��ƲL*;�5I��D�(ȵN&���nM�pn�4�J�ަ[v6E1@����i�����x�$��`I̼N�W�wh�_�ɞV=�>�l�e@	G@��mt+�?8�O)@�������S��an:������`4IU�֕��4�n{�9�|�)T����f9�Jђ]R��$X
nF���aq���a��t���c�#"�Sӿ����ݙ\�����a��h�qH(n�s��5w�>�$6�n�_�LR3	�Uv%��E�l0�wd-nUVƄ):�������]��FϪ_m�^D5�*���rBa{6g�췰�J���J���<�
,��FX3�h��L�z��q�d~a~��\b���_�D��m\�݃��k�ej�B*\�}6�}lQ|H��QP�������A�Jˡ��(��@��[���&��Ǩo3S|t�0bL w��c8G�]��C-�І��Q'�bۛ-�c��/pQQ}N�B3�g�+�d������j:7��0��㠤����5}�-�z�.=�;��ۘ��D���~`wx�K|�uY$?j����p/yh0PH:� :����M$4�%������d5 �Nb�zf Q��rD�C��#�3J7��0��A"�C��,%�f�H��/?�"
5T\�#Vo^X��U�P7M�d�����]�h�3wy�i/F���m΅��ۄ�Q����tx��,��R�q֖Q]�G�?7���@���2Ơڕ�~,*�>"��=�h��<�����~: ��V�`2Ҿ�]��9��4y�'�:�9<Gޞ�L�{9�G`R��.���>�x�x���No�z��p_��l����޻Ŷ;�?��dh1hQI��u��[;���ˈ�W��͊Cn��)E���q?��ݷ�U9މ�\
�v�'/�)p�|������H)�C��m����|�~�3kJ����y���V��1����ڊ\������|T���4���fM)��tK|wCK�"_	��n�C�=��[� ����%��j��	������y��