-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
KWuLcWHhFJ1CMVhXShILIkYYhqeNGs0SWe+HQRSgNfAtOgRqJM+hk60iQJfG4g9g3aN1O0FGJs+e
JQqtk3yM5O2feVNwudzorVsbStFGx2y/GU4OQk3g3BjcEdm9j0Ybwjfnlv6eHYX+qgJY+VPP76TO
Q4Qp2G4yRm0Y/K2FGgi8COK+XgybYj5SYA0Nh1s+DT2cIAW181BG3VcR+3jlvcaj600M+QCVXppN
oyZiKS1Km9CjYpnAJkxNNBb1HtxPdVRr7EAeYk/LbJUJPQxz4Tr7SLA7aaiVm7Ec+RJ600iaFW0/
ACzmEzDbu3at2nx3YcXatZwRRN+duQ+BarPmsg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3344)
`protect data_block
B02qZIEILS8GK394DtH6tXU1DHgxOs3+dpb1iKeXrJKFU8AEZx9m7O8pD5IljcaCdxHK/dGo9EIY
sxdHp6X/fho5u73oRjqBV4uGP5bavVO8Vp2Z32mA9sPWvG44d/JfUw3FHAibbzbtB9SKqrgM9F3x
D8RrsR3d2MFjENDTwe9WVhD3QyO+KQyUNpKsj6tM4lKOqG/Lj3sSzCLGeyC4Y+Cv28fl7bPYDrm8
O3qPB9HzyZpbKYDLSHMrz8ZCFHQFKVSGYJR16hhy6P5jDum49WowNbIEtRy+xm4Ts0VZtA9x/16k
gtPgie+iPbBJPseue8SPOnbQClCBUnYzfbJmn8saiddlT4XwFlENJmOFm7BsRHkMKGW3TiZ57rM+
xQX4+wtC0ucSOhHVdnFcocNeNyYpw7cClp22ih6pOcIVqYakaMBeUDRHOomasuPoJl6c46kM7gky
kVnWgH6CusQbksMwB8yktET7ICEzbU2dxikoQRWlYlVPfO4j46Fu6AJFCQELN4mkWDssoMmGb3Lw
ZKZZgbJuD/BtNqUyeFms5HTeOu1uU9ffO89yctyB55VWpnEBh+LJn0ZCuyPAZWV/bDKPpJn0oe8x
adtfduA2nfeg8tN74XjYRjPHQT5X96z4nwSpFsBXcy64EEpemsjFa8MSQ8NirGQAsvK/doLx8jfY
yXo66uRgT5OoCplSFqpsJd+gg3n77BNDJ70OHbuvBfehsJpcQYCrA+l/BPFGYh3P3OoovU6xhPJX
rBeZRYfayti5p19KAUppXGQsX01OPQMjd8dvidR0wyhqY6OhVWi1JRqSfEBefdJ1m2f7204jt92d
hHuo7V//hXalRrPxvAiUdOBh3VJtgrlbK174VozkMrT8SjBmOqZPj9TlwTOOSk5yNLlbRnmEmsa3
djf6L/v4sU++9JCaaYmZ8rxqYpCXbYrR8H2Ez73yQ6siQUAU5XfoJtOVycc2VTfymuxgu7si/ted
HCzheR6vioU7eUWeu3Vv/2iUAVbmPnT05aM2Si8uantgQ4URDi8ui33v+yp9fsvpr9Ewv2wBMT/3
GHz8f/FAHCjPW0fawELzjiiAwowGf8tD2ZOLqVVkbqY/mymviP5Z1UyZXFVulGwwtADIxJQIb1v/
UNx3bXlE9w5bLcTOCVO2qyCon7TqLbSn3aQNLxPJDrRox+LybBh4kg0ONKZzUysReH07TJawRigw
4FWtZZA5NYG+8H2jjPkXe+QgI0P7shjj+dMc1vfP8OC5Gcy9Qb4M0igkLzPsohFlpIY/FEJeB0ak
VoKplUSF6uGZpuhVCUMmVcuna02hl+Pi7bbvp7qFm31NPIO02ANDPtYoYGkEGbC/rlIXbjjOJRQ4
9jXhpo0d3trxkM8Q33hEeX9xIQz7+cA7MbnBaWqbL2cp1JUTmVIFCykoegQMiVDx0WpWKrFajiGB
LLGO+qWc9qA1EsWuduglgZxDPdl5vAPtDl4yYkCBzZlnmtyKZp/BDHizcAuwTL/gNl19F810PX3P
ncLRPRAMr2SUQg1bJShy0HNxx0jed4goAngYobMp5fW+MvcEdALCUg5kx2YxcoflbTPEiX0J3QEr
h+XsV0FUDibFrn+90+QHMI+p99HE3m+a27sv+0FxOZHnDY4l8bxwCCtJvpcy0bfNViCsgwAztt2l
PLX0bFwRPlSVMItNVr/+sQ34kgT+R4FeBroZTOG2eIBSRvS7YWB96ixsQQL4/fpaGKy/vH+mBjtb
8dWIth/AglSvTE0wuflXH38YR7jm69PGidJhCoHQanRBIfdM2cb6G5DolQh37nK4NXGuMrX2Vv7t
TE7856Qy8SCl3d6I1tFx571lvbf0oIquRTjtCr0kQujVESxEWsUkB81M1LFlp1Uo/9pPcCI3gugW
0sGv7gz7XpZSAcu5N9bh8KWymNn3tt55tTEs9jy1ZV47w0mx3NuYApDU/ljlVsSBXToAnkuBbKqd
CyD2C6Bh6yLYZ0LLa08+95hweRCHWG/Hb92aYONUJMONiqKWyfkTj3vCMQFUumkw22ThG6NKP5+7
txTS3l2Ir+rSUYmQuJetGcaWFEQd9tEGDyAyNAQXM+LYcg+AdWxdCBJZUIZ46gbSTUnWnyOQhRK+
P+AzgXJ8iRGwadNv5pm0wpBNR+JgijarlR0NTseb0+BbK/rZqYJzRMMtdDDybxtvVfgzzNzX4fZw
31JUvuvRXjTtKfPNwaj9SFYN/ZjELgNiuuJlGj4ijRM9F8Fpjn2ey3YkLZbdo31oNYfIYjCX5s01
3HzHyiTnGDd6FdSgugU8KRh7HF2VjzBDBMvEnFsL3VLakjyQ1vALOp5gdQ9Q3mV8ViwLQjYIW7hP
6vz3kmDoVkic3FayNYOSdZVAWRr+dTGtc+vvk7r9Cr0LVtaZ31Vz1obC5ZcACIE4gzyGqV9TPXjl
fY7t34YSdmWLo/Qx9L/Ond6q0HEPksj9+Dx+YebSokL4hF+eHbYkAI7CFiuC7l0HCR7E5yswpVxv
eBgrl42cRVX62pMlCKMKyKU0W/0qlbj9aL2PKZ6TKe8DFkhNmvMFPqtxKJ69GyLGot9sshbuXNDm
G7TTA2ZEY6BhdtExZ5eryA8yAoUf/pz0ZtTkgbyjnd41HYbdZ7WRpBPLWKdT7P/VIib3rVWebCbu
tlqWdQfcVOPm104pG/VZlsPfPf65yPaifQ3jc/+ulw6QCPtlDEnaDd3hNZy9AQG3IIeWOSqRhqKr
1shG0TmxSbu/hWItWLC3r89rBJHlmpNWawAb15YYV6Cc3OOffbFAmeAN2IFmQ4VWyvjfazVHwVRI
nmOz/HQl88v/EtOpp4W8Z5/6E/TQK0ZDWYfAi3bGyyi6xNkLGOZYGbP4jpjCip5QxLvp06EkDMwL
kZs03yd+Vau5wBE5bhNY50OU8XTaxKD3kfD5YEcH1JwPvtRJsyvTRceRMiCUqNU1bnukPQRyvi5t
U3SmWTaINHGA660vIT/h2O/DxL3L0HPfjvJYAPbg/UnEFfRayEJv+zB8ZgxavCl5Z26vVfc7MD08
0QVLkG4q+VlJ21ezTLIm1/E34sc3jedVJpIPyhV9OEC2XZRUVS9DAxbSp+vzMSuu4y4s3YS1qpx7
rdBr/c+3oJAzw6VTG9HWZTPd6mzAOxrllXymwV3glmSvJ5F9JSZTX+6N15eB/flrWvHsCytsDbFz
aoB1+HgNTKPQmH46hKfsdlp9OQWCaNv335KqzohQJlFTzLmPWoFlWAHUidQ821EqF8FpEflGR07G
eqpAOMv1peFdgNzIJkh4otSyLF6vKC6wUZ1d7bSWYCYAxb+KJePMx/mla8P8HIKLa0GIh0v/YhRC
sMXW+TkbbsqR51m0ze/Fq1GVtwv/+12tqvSb/eiqcjs47s3kMX4C6YZVcCtG/OPTGUTTQX8hfNGE
Tbn21XCfKYqkewv61nsJeRLUAoQffxPFaCeW+OB7V9ABD//18bbERrXx/nFJY2+qUBp7HFE8d6Br
Yh/KwwRMyQurXqC3IwDSMynHQMavTYr6QsGOSSskwC2gHtzlmQ4q4R3YF13kDU7riv17nuon1XT8
DSHPBkuDccbwaOfkK9RUT9IT72lfqt72HfeLUddHZGZ0DEwKFIx5W8L7bCD6xiaKJHZE5aNzJKSQ
pYKZ7KJ7VP/xT9ytBEWxZyzTtE5fM7J+BhN2Saf95l+HKZYBNQB1vesFJS5QiWCo4tYNKoadyHtz
fnk6axr9W6jvi16yN+vjtXFK2Xy6lwwIeDl55gaDwGiF2/PdZvWmkhePVBx5rC2iw6d/UhVM+jm8
UcInaQsmZXbaerWDYdPACnEkSaYlr4DzwyTwQPA+qbb+0bD5WhfLiddygdaLvteFG5OwspRrvb7f
MQpLeBbXaSUfBlC+KHHNfqCRp0BTMJy7WYp2Ip1Xbgosv+bpfpk3yEU6ZOUet+I+1tKxlsUhQBCg
YqldFz3zeulaB3pcMfoSgDFVPdguLvtNtmDAwicb8fV3I1ScTVfsjfepUwoLeDuAGvzIxFx43fI6
fiotnfiVBx12KVrvbB6cw41cGyZsSU6GYPZ4PPWQvpvPg2ZqOW/703hv2Fla4/BaAsHZ8sXG1WUR
LPqQE7uUs1P3RadIS76xZ7RV/NxxuOoNi4+9ZZtnatHe8vCLqBqLyePj15JeBb7kM6o2uliVdzEU
CsD/3Drpmai/scCn7lQZQTWZ/SRbVSXfYVSLBNWK4FpKptyEi/EgdrjUO4P9ikZJIA9jdjsgmBQv
NT4F9FeDHjUHX7FfEBzmk/+5q7t5kiMo3899RA2O8sVk8QpTXUD0KACMzh9AozgTt4OVXbaIptj/
gwwKnGN9v/BrYmbq3t04yRd6j/5/t2FBb9uGymEJ7vSivpJA8ocwBa4zJCb/5igH9I/OCM5ejWqX
5yIwigk1B3F8CCB4PhpIpwUq/hkirS5Bha2gyzny0Jjf68lnpo8=
`protect end_protected
