��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[<.[tӒÓgx���)1��i+�K�SY���'o�yM6�`kNX�
���{A����R��%�=4��o�2�ИD��ȓ�}��t�z�-7yD���)C��<�f��qF����e��I���8�	v��(��z��{��WN�'Z��w��&΁�R�~�%��Hp����U�/R+f>"rE�;a�=�_��k��L���GEnfF�B�y�1/3��ro���1"��� Q6�B�e��*|&�<�%�7o��(f�m��_��Fr��;*��y���ڪ�f���$���%�q�K��4>�>j���Y�#馞v;C�+�W���S�-�H��/��B�U�ejpn��N����͙ҧ �X�|`�w����jl0��#�䒛������>0^�ҧ�����Yg�77;�M���]M�lbrs�@�6װ��^���W�'_��� ێ(�IZI,���n�4�֥����'��{8@�:i1��m�=yl(\x��1aw#�~� �(ŷ�RVy��,�A���o:���~�?%W�wT}(V����+�ʶ@I��S��Iű����@
�=Ev;:��z���$FEZj�Ja��ȱ�z6<��1�uxd���)��SeI\b:��d���ۗ�6����2tə�e��i� a���<"�h��$}�)S�NO�1kð��v[!�,�ÃRy�OG?`Zeݮ�^���Y9��l,���H��+���O�B�L�UiQ����nh������̖�'�?C�$�)�^`W���bI�蕻~Y^0
t{�*-@�CT*h� [�����F(�\2E����F�G�9z�8Ã2ֿ�{���
���٠�t0�\��͋�qgW9���O�ِ?��t�8-���xȾ";|�-]���	�}o{,����a���a������F�Fɴ6z Vڻ�Jz���(T���j;�2��}j�6ˬ���G�#7�5�S��<�����o����� ���9V��<"c��)����t�|�R�v�3�?%l�}�t ���r6�H�{���4���<�¸AL-f��Wkj�C���G���BZQ�I��S�?-��u�Y�ђ+�� tpi ZK�y;����fW�����}�4�V�H���I޵��]��l����`PZ8z|͚Kam�?Ȟ�P ����i�����·��xq�h�����~J�z��K�_\�B	�ؘ�8�rS���#"S�E�Ia�enB2��[M���R��T�����7���b�,�B����
�B�.��,X'���aɦfY�B��Q��:Z�!�]i��D�zH\1S �;�*����%%C��4}�ԯ��9,�5<^����	#���Xl9��Jի��0$E�O�>G�[�A��f7�=p��w�Yv�=�.�;�Q[6	2�%��Ȍ2y�$��K�v���ʉZ/EZ=+D3%�%KH�� bU^oQ�!�+|N����~Eƛ���Ϊ�
Y���W~��q��i�G9^-]�`C57��D�J�P@r�`�Rܗ�G�.į"D���᝿��~OkH�ǌR���,��:�X��Q��)��?Y��7�Xib2�$y* ��<�D��{���Q,��㟃�ddI�0%	mGY�L�umi�)ڔw��}(�ݰh׭��K�ŕ�P��g������V�~}j�K���_��9+�+XZ����r��!��׾�Uܥ�g�_�G.l�J���v	�U�'d��u>NVO�C�j�q��h��L��U2w�S-��<2���h�RH�nK�s��y��n�������T�ޝH	����b�H��I˝S Hɟ��Ll�g�~s��i"�ǲ��rbD��@�XYĪN�{�@uo��1�{y'�k]�^���wM�eh�w����}]T�ٙG^�P��BP)�q��J�������DN�b�
e͕tpєFK9$#��W�J�j���ľ	T=Q�>�xƸ�����6�9�I���hYG�ϣ�h�b��	�Ϯ�#p~��+�cAg\)+�gSQ�J��KO���^��%�[?a���^�TŹ�t_����+���z35}dI�Ŭ��y��b���͒�,)\n���iS���2c/�&�f_�g��j��6��J����ժ5��8B�u����֍��fs�Sݽ�	�l#-|�>$�ж����h]uESu�q��;�_栆L� ���8*�y�×K��	-��kI&÷��?��1r���"��x��-|��G��'��*�L�r �����R��*�ң50�Jsj��~�JMZ��P�Ʒ�Hxi_ZF3p~*Թф@��Ѓ��K)�ձ���!D�٢*}����Ea���UpJzi�R�2��<�ODȆ�H�D�������H��R�Ǩ� ��#S��pr|le�%�	0���"|@����k*�m�1"��	s��-z��=�Ɯ)����tY��ri�(�M��d�����L&�i����5��ܽ�J���ڧv�S�7a�Q�3�Em��Q �e����+����b"rUՒҵ:��O�材t8\�s!_X�	��&')k��^Bm(��B{L3=[��������[��݋��{~_	�Py�"+C��׬��;V+�7�k�ꖾ�V]L���v�)�w�-��>ʗ�Ŭ�ڨ�ɩ�D�ٿ���r�$Wi�8���1�P�i�&HQ'c�Dmt�m� ��_�;r�=�;�����f�J���H�����D3�zE��&��W��zI�����,m��P�D�e'r�ܪ��mm�T؝	���w�~�?��TЎ���Kȥ��-�NV�׫o�V�㪰�(��@��}$3`�Ϟ�C��Cq��i�>Y�M�Y�	ò���j~���k��ˎ����>" ������N�����ɭ ���+C�z ��%�N���o@?����q��f���e��G_�HY�H�6�:X�Re�;Y�8�1�8���9~~Q��a����&p\�[a�</ P�^i�y�(�ʬs�h�=)��Y�c��߮���@d���o����ê���`�Vzﴪ��� `�?��J��C���B���L���ͣ�=MG�ߒ�r>���	�E\������F�2���%�AeW�����^=�4�(�����8������B�5�h�Fl�4��Z?�o�ˈ����/2A���4�Q������}2��A���MWV����vڍ؅�U�<��P�k��g1�0]q��kw���~�C�t?�_'HPۧدܳ�T��\jn�?B���О����헫�`�T弝�����\	���jC���UT��#�~���䔈�� Ý��g��ʺ'�X�o��V��!p6��/i�D=���J�YC�bNR����t�zY�=��� z���`����'�މUA"�Q&Y�gYc�H|��-h��D�"�@mό}���c�7�a��ܵ��&�)�ݹ�M���4��<����h���\�z`��NP�x���"���2C�u��Zbln�,�R-<�4fy�IDؿ4^ۨ�N�#������Ý�܂�$ك)���Ry>��Y��*����Ī���%�VPF�e��o���7���E�?��`/��=��e�c��(��>K^���s��'IY�N����&��f���R�@�h<����$�VqfOOE��;����lAKYm��=�o�g�CL�wVU13���}Cd+It�}�n�5�v���[�SІ%��~-9o��o5��=q�����U��:�ep�Nn�|�\���$�?:�1�����m[�(0�4;	2�.L7���j����_�������%��g�)S"f�O0��"ۊ���R�t�xOd)�J�[�z���ZLPM(�h$=v�����v�0Ka	�����6���&�U@R��ZR��kt^]%*�Q̆��Eh�J`@���5�}0�����>
��d�5�!�Rh�gJt��S~�	�zm�Ip�Z��n��V!�W#�J�t¡�s#�� a[�m��X�g{1�	7s-�;�(G�I�U�%�~��.����G����,����DI�E 9����LKֻ�FC�^�J��ƅ��u�~G5^���D��B@_'Ŝ����}"�x;��xG΅Q^�޷��q����*8��m������6p\��Z�(v�	�{��C���`g��t3�ʹWK��\.��U&~�%�O[S�8��U�p��ھ([��Rn�WyrV��J� `��BZL����(�<�I'�#�:+��<W��%.@�l�$�����t�7���r����r�%IOg��]�q��Y6��t��y��!�̘�x1�(��chb����4p���[�b9��h���t�[��ﲶ@}«X1!u1�7�#J��I<��h�5�%:�썤\j���X��<�Q�8d?��^��N��ksC�A���p�j!��Z*Z�>���6�dnQ���߆"�`�p^
$���O�*5�&`[�!)�A��3�;���b�=��"�J��vaˉ�%	�=�x�<=�:��1�ػD<�Ai���t�q�Ca5�cg-��r%� ��lNKD��G�w4�Q.
wYl#��R_�4艶��Z- ���J�o2��Tw��OSf��R^)'������ןk�e�Xj����͚o�48���������*Y���i�l�䢟�p�K�OS2��|'�}�/�37���i;"O]X��[��k��v5�$�*)���]ҳ�q�bw��DZ�ѩ��|[	�غA.pb��k1o��*dN��l����9we� /��k^m��`\H\�jS8�/*0R}غ��$q��T-2�#�liq��Y�=[��	:���'�X-t�:}3��q�Dn&"���a������v�|�|��+�U�z��l��U�ΓJ3��=@}��*Dl����v��g
�TB��¯�I�����A��h�G����񦈹%2A%��]��C�o���|�ƀ>R< ����۶'�
���V��Gg~��Ԉ3���D
x<�%m2���`��x񪣲?�V%��2��)a.�֬K��\�ڹM0�=^!r�ꀞ3���TF�Y�9Q_�N�:�2�x^B��j���� }����x�u�1���[�y��?=x�N�&Rvx��<'}Ҵ��rr;�ռ��Y�uoV��L� �B��&4*�LCVR$���h���lĀ(!�ҏ;�Ȯ���}KO��\�����\�;��*GZQu]�p�gp�x���?��)�HA�=�k��c�/=
T�J>�����S�k�s	]�� ry�U�"�̇�qܙ��z���H�w�y�!N; �(��d�_3EI����M0��A�b>��7�L�y��qLJ��	�Or�����Z�}�np��}0m6r�I%��5H��,U�z_#�}��~�b>��j��
�X��c��W,�ݳ�X���P�(��|㇐�,JN�F���iJ�F(&HF$,+�6V�ʗ�L�js��.2�v� ���BEر��U�M�-H��TY�6zf�i(|��`�M���o��'t��TXU*�Q��b��k�����a{:�	��^ �;�Ƒij�J5d��������5��
F������yUJa�kT��n����{tqQ��,SSޕ��ȑ���p`��kzn9�S�=�E߲�攑�v�=Q��9�L>v{��Kӊ)Yn�Đ�TӢ�0Ɣ�j�@@3[����G���N���`G}�t�FcV2p���/���24r�#�)�j����"O�$�+V�,��Aǂ��;s���}�ٕ��(�;���3π�473�`0��ZѸ'�k�(y���_+�a�#��:K-2��ƞ3��؝Z��4tc��	N LF�o�E��d�i�i�ӑ��vcג�_�vs��*&
_�BZ^������O��혴��q1��iW.����� ��Z��cU��tu��B����9��1�Nw���
�j"r��#�"f��*�s���{��s�ټ~�]�
��b�%jc��<�A�~0;'���H�r�87m�mۣ0���F�=$�q��Cz+�{j�`�'��8�m�li��7��Yjq�46{���!44��g�*�b̅`�ǯW�-�=c:x�-y"��D	�$إ?0xhl���������ݔg�0w�S��q�O.��RC'���Ű@�bz.H��KU����
yJ���fq�p3���ˑ�F��>�5v�^��{vye��Fo_�V70I��8
7b.	���B�_��+n9���Q����(�ê����%�=F0�c"JZ�wɆ+����������c2�8�$Ü'�^eM�t�M��s������UF[���[E}�8�ݝ���,�g2��Z�]tY��*��O��ϊb^�C�/�bHu��X�jq��M	�G\e��}iG�2V�U��i� ��5'}V�/bJ��o[��A�I�<���5)�C9"�
*��}\����W����k�5a���l:D��n�<%� "h?A\��(,W�{�=s
>��?|w�#h.q� ��p�JO���#!L�a+Ot�|���Sͻ���j����PR�³ć�����x?(_Qh��,p2xG�眬�q�u�S����*�r�v!_w8&Sݼ�0�K±�����9�/�!�TH���[շ�`)P�j��;sQۣe!�=�4�������c��d���c�/���{y��{tf7�v[�719��Kl�ײ�#I"���V:9n�եL�O�k`��`�����^�@C9L�.n�r�f�e��q�#@O��vc�e�l� m4`�\3�sZ�L�������4.Ķ���y�X��Q*g�t&*��T��oR�߆e����ؤI�1�}�6�,)C_��n��Ec��m]�L������(�������)*-E���xU"
2n��v_��(Sv�XW�����󰇔�
���T5���׆H�2���)gP] MP���3w���֔�������#Ӡ�u�(���J�H���S�Vv	UE�g{Q�6�d��U��B����W%H�(�7x���ȡD���$�c�Ƣ�������³����8���+��\E��.0�E4�@�w�u� ls��l%�*�MݸP��?XDAҚg��|��`��,)4x��Yo����1�|�{�L�#�K���F.��A�ڴak��B�p8���]��|�c9������4���I�)B�5Je�'{L4�o5^��u��y,��nە=�(�\�J��	��!�e�R��C�.�x߄6�ͳ'џۼ���n��%K"O�@n��N*q��� �������ጽ<��U�>�;3���&�bp�.�M�C���������8���V���N�a�鬙�3p���]��X�q�`7	��<��K��; �Y��ga�#�*�H)Rȹ�Af%�}����Wpު�ف�U���)��}\8ض.��K�E��]�qW՛�>�v���4�l�!�G~��&�p�F9N��s��>�Dj��i5�Ë(ʥ�p]�\��O����vQlv�x ���q�.������m���cS!��$wC�X9x�si$�[�-�� f}�g?H�KH~~��̂.h�]e�$a��:�Á#q~pI�Jt��_рڕ�e�;�d�*�1���u>�t�T�6��	�D^�I�8ˉߒ[<}��!�\].Iu�!n��ي!"h���*	ò
c�z��7�I�����+���u���>j�eG�x��B���i2���]9jS?6 W�<����O��3Hݹ��x�q0�3��ˇ����!;Q����Oީr�m��_���$�n�TF�;g���]!��b�\|���p�@L�� V��0�%�N͕���Q����l�A�LƜ#�}c9���y�\�~q��a-�W��Un�-X�������d#-����C7��Ųh���-�V&���3�aK�#kgxʸ|B4��������n�]�l}�VgvS ��'Xh6���qd׭s�+8��K�Q$n%�v&��l��Cq��i�2������I�ަ/6�6�����kg	bK0�fq�v�"�$����;�Q��fC�-��Z���gFΛS7'�~�^�9zP�P����>�VO"	��p�co�U�O���4ƞH�6� [��	�rߘphH*�[����ג�z�Uy�kO9B�1.���� �ؔ�.;o�N�x U���J�s;�	��1J4%�<���~įr�S=cՓ�SL���h������BB�r3Iѷm�L�VH��9�O�y"�f��L����b��ds���o���nȥ�c���g��`��tN����g��`�:����(�H�k��� >��ѷ�A�c���k�=x+ғ��dB0�Y��HC&7�14���Z�`��wQ��nFS�eo�����͖��D�U3�+~�w:p,���gu�M�Ȥ�������A5� i�5��u����Y_��D��
�h�҂dH�L�l$���]�?6�O�V�1P}
�Ґuk�����~i4��w's���fNm��m�9MZuy� s&���M��J�?{XP�M����_2ϵ�\�Cݸ<�r���JTcT)L(����������7Ozt��H�X�7I΅Z�]ysG������)�e�P�rߔ�D���:�m��F��|��i����5�S�?���/#T����o;������Ͷ1ew��K�DY&�	AC��-� �f#�a��c� G�ީ��

����ib�B[o���3<¿�yF�1�]�ko�~��q���|h��QL���p�J�ZM��s���y�
=�?.�G�*�o-V=������9e�6x����dl$<^A˓�sR�s�`{���^9m ^0�|��ڒ����B��|��>o�47��y�85�
�}D���<��g�
�~d�?/+�Я��g��ν.G��+�ڣ��vn�L#�G���[an�E��i6'�%��@�處ŨOMDK3�H<w��R������g�\�I}1
�=l��IzӬ!�7�`	x�#\ꥢ�鬶��9@�f-Ʀ|�[��q�_r�V���Uj�S���� �I��|�4��,
N���u~!Gm��U��ۀ@�E����������ڈSfr�Ѿ�;g��9�/�U��3G�;��.2�m�����6~?�-�����}M��c5��}?׃wk�<��Z�aI��W3�r�M��Є����{ϗ}fk���X��{]0���8q���a_I�&�1 C�/z����mf�Oج��}@������S`�{����դ�I�=��t�懲B|�~8:�t�g�H�ض$�A�@[�TUzڟH�ms{�!ߕΈ�֬����1emE�	�n�;J���׭i�#�@N�K��?8��_jT��ou�R	��zd����yGE}�2�P���S^���ףJ�s�*