��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR���[{�T���CK��TC,���:�
&��d!��]9�'D`�"9 S%�aQ�`!�6������V�W�l�a锦E(�\gC�slu�4U5=1�N�m��l�9ў��P���B�@+yg��=�}|֦���ָJ�br(4-b��!�� �1^�l��pL��)3S�(1#&nJRę`C���Ų�����B3��^"����I�FU��؂5
r^�QZN� Paѿx/$�a�N��D.�Y����I���GHYj�ݯ"r��
�WOD>��k9��0�Q+�&>o�2nA�U�)+!��&t����y)�[ţM2�e_��m��`V��"�ja&lv�oF��Ζ��~&�����Ԩ%y�Kt�g�/I^�I����_"Z��T�Z1\%6��u���#�������ω��ݪ��k��@����?}�z���a'��3���|G�z�����c��l���E�	�dUp��+	M�@?/��w\�O�~r���s��Lu5�����o� �ۦV��c�H�BS�Z?]���+0��<��*W��"�M�ik�����~`��3�"�a;e:@;f!&��QW�2��6�Rz6���x�R@2�j (�ê��J�ҥ'r���DZf�w���o����nZD�A��Y$]�1�/QF�o$����O4���.���q�>�	���
:��IY�1��B��a��Ս~���",�:kZx���f�R�K3T.�$�6��f�fyh�(D��]�n��n)���M|؃h`���mjٿ�e=}��B��h�60���`����@�|���/��,��y�T�� 8z�0_	�y�E��1����$�����ǉ��B��F�{�<'�,Έ���ܜS��rj�x��ȓ��]�$'_uً�/(?�4���1vP�S4h��R���޳VA�K�z�N������K/'�ͮ�ϐ-�������[���K ��>��=4�e��pᛓN�>Y�J������jYzQL�K���*�mB��/�\��yr�e���N
y8�Z��D`Z(�$F�Qj�w���7w���6e��@Φ�Q|-L���j܏�U�S����'bFS�d8��ߛ�j��U��Q`)D��L�(�䆍4��A�(�{z_��|��C�;��o�7f�c���:��]����I���"� r"��$wʟ~ڴ�Љ�8u�������4!�ņz cC]�(��_����
 �kJ k핅J�f�87n���(�r�z�%���h�ΈۘI5���qB��r��/���eK�:�>���+�I�?[GڱpGb������I3B<1������K�LAh��D.`i,A]��&[�֒�㙁+��1?&�0��@��;�֘���E:�%v���� W�[���#^[��N�:��A:l��wd�Mc��=��6��	-`"���ЧO�Ӷ��]u�X�"��˲�8��Kҏ��>B����ar��[Oɟ�X�r�k�}����}r��J�8ېu����쓓##�����R�KlC��+�����b���	�z����S�ح��{Ǭ����w��*/`3V���@6d�Ѷt�ƞ��cJ/�j����7�[���]rPl�A�Z���5�?v�e�|���A�Sҝ��
�PB)	�?�ح�=���OE�(g������'��%�Z4yZ��6w�JSP��h��b��Q��Q�)�HJ�p�
Z��<����V)gvX��(u��h��q\�NVKծ�A�N�CW�+�:j�h�*wFfa.f`�@e��.F(Sp��ͨ�q���·k1�	�y��^���	,�����%�ҷePǨJ/�67�;�+'�dk�}#8Ѥ���ym�{( 3�F&9��ڗmU�W��ím�\9�������!��
$��
�UzG�"��&Ѱ��3����x�aPA��s�֕�n�4>V$��zÚH������s�dJR���;\GE��r�=$�ت��ڶ^�E^V�����ݣ9ܘ�9��SQ9t���u;�neav�F���t�4ׯ]����ς�tHKc�!�
ʥ�����p�3Y�"�	��w��gO�h���m��N`8,r��dq3~ڽ��6V��	�@c�{��@#�j��\��T�S���vǧ�]�H�p��O���;�zȴ<���z�'-8�^q�֤|��r�@�o��>u,�mN~�4$؀����f��|�/��BB�5�U�c�p*sC���
sh�%\	�R3m.�ϟ�i�}_X!�R�uaJ��8ġ� �;)�6�s�h�/~sdj�ڶ{����ӈ:��d��k\.U���&��vK���]ՉqIyѓj�FFc��)
���٠q����V�4 Iz��2ʅ����$�$��}��)�y�AV_��IS\e�xf���V}`�l���v���s�Ċ
��&�8&3��a��>��op4h
ɪi�?pb��{,-�{E�M}�ѬQ��"�΢[R�a8-n����G�(*p���^S�#m���r�A��)���U�*YZ�����v�+���&$��x�6���P?���s�rz? �by\Qf���e#ۭ�F߷�#�5_Kȱ��*Y��q a�?��]_�ώ*�����w��R�9�?�׶nZ�zB������^B�5m2#���>
Te�0w�����!��9ӄ�i.��C�@k�d2b����g���2e�OM�FTko��(3>n�����6�r�;���yG0����c������uźɺlZP	��!�5i��$���W)L�dY<�}��&��f6[�!3#K�(�{$�������k�M4M����J��!~���䄨���ɧ��$�b-�X֊FC��sޚd�GK�&Y �gB'�_;-8d�@%���nd��C��ɡM:3����L�Uf���2a����#>�z�/g�~�����u���"�{3=js��3�ַH[���`��Ѿ��(-�V�`�����a�T>��LԴ0��o#Iv�r��f0X;�����N���k6�o��jፚ?V9�"�e��K͐���>p����l�Զ�:8h��a�<6ӎǠ8#�6���pf��A� c���Ey*�$@7C��?El;��PM�� �^�L�t�c���5M�%ݧq��4(���*��%���@�ȋ�Nu�9���.ǉ2,��\�]�	|VYv�z?d�KM4�_�f쑵K�q]4,\�fPȮ�H��W �-�ܲ)����$MYIO�N�`U��T%��K��eS�Z2�mx֖�m/�ϑ����E�
-�z޿�9��p��Y�C�r-�h�7ȸ.]���R���x��N�Ȍ�c���K��͋P� I�[���١�n �?������ ���z�C v���}�Ie�:Zȸ�M�F�jo�'0_dw��b�C�dh������'�jxuCI�6�Aj���gn�ΎA�k�C\�t�[���=m%X7J�>y�O`�"s�yü�������������3����*)̒��.�oڃR�[Hѕ��.����L7��V��6z7&��Ty��7/�,'��O�v!G.u�x}o�hz@D���nJ6��7�4�<V�G�^a����\^�aYI���?
�䫪��b���ݬ�Vm�&���8�w�S�L1�JZ��QJ�`�wc�SPZ�:�ƴ'���y?J�����3���� Ű�b�؏�8x�� {�%>�Y&�Z�#ʆ|a�o:�|�J�ԅ�U�g_+�
4���.ճ��j8!�����d�1�`a._\�Fu9��`K�P�Y4CW�S<�`;Hdy�7B�*��-���#�W�F��TU#j���18Q��`�� @�<��a���U�h��f�q��ۀ�A�{������H9��6�k����p�,�& pe��,s�^�ir�`;n��(�Bwߢ��bG*W�K��m=z��f��]n���1í��RM�����p>:
����bo�<���zc�X���^W�-K4�r�1v�c�>y�&�杳�+)�{��SH����53�^Z�<���Ѓ��W�_�J�#�Y��в���y�+��=p�Y*:��F�ޛ�V'�{�2�����F�����j�����oG{sѽ�]�w�:�J2Q1�o��H+=9�i0D|\���s���@���X���ka��E����Zm�����m
g��z�K���o�E:�#�=��>�X�4��9|����Z�W�7v���/x�����/J.��@����K�&Yޠ�w����2p	���� ��H���P]����H��ݐ�"��E*��L�u#��(�֓�5�M�vm��Ò���:p�����i��vz(ȑ�(=��A��i�s|���Ȣu��oȤ���6���hم��6@��� ����׬+@�O3pd ���G��+����B~a����X5o�M�_~�É]$��^�άM?0&�H��̚�ab��$2��fe-�JIO�|�EG���;�^���qZ^�vyب/�m���W�.�����G�\#���e0��uȽ*,�*��8w�=ݦ@=VAd��1�C��G6����G�ȯ��jU+M��> 9���Z�=#�]J���:�U	�^$��<����S�l�b�t�^@��^ϨU�����-.�"�1�B�,�����o������ǋ�3�}�$�6��#+�P��/�DU�~u�`���z�����Fp[ݫ r3�,�_��ӫ��l#���K���|(����p���E��L�����x���	����7�o_�n���eZD���x�>Z�d$�O�Jꞵ Zj�u���eF��v�E[��ͩ ��n �40`be�]�4^PWj��Y��y�>仌��=w��gg)�kw���;�4
����6{�߉/&~k`EL"�"�nYTeJ��1�ҵ���V�&�ՠϒ����uf*�u"�Ɛ1����������[��v-b��c�K؟��59�8�h�&�0�Q��"a��X5{G�i�-�lK��ۓ�����
�הU�(���5�5R�2"�JeC��_qq��#gν�J)ޥzL�9��t�v�g�V�Ƀ�W�\���˵�|�6Φ���{�9�uݬ:���xkv8�6���.�v�_&�6�P������bU8�������E���?���v���-����}Rʅ��sX8�¯��=��SmT�v�شu��F��xG琵8�� N��4 �� ��5��S���|=+ɝ��yAɶa3kt^��s�~��պs�sx@c7��)������{r��Yz2a��o�����
L�`�F�w��{=���*-wN�~�CQ������tz�I#'�CCwZ47|v>����X��"�5���s�F.�J~H���xq���uN c���/>���93E����TU�ʪa�}��m��K��g|HЛy��~{�+<Of�]4-h ���t��@�*cv��,�|;�B��HRt�I�5"��++�h~��lj/�h���aB߅�'�D�Kr�>���sΐ��
�Jn�7�!h?4]=�}U��ܿ��}�X4�1"����Υ����a�a��"�E��֟P��O�XƜ}2�e�āo,�T���#&-���xU)������`iR��D��eS(˱�WV[�����5�UxX�� ��ױ�z�uNu�:Dj����Ms�%d�I�k��ޘ`u��T�;߈"�*���^��QD�@��!�)�=xS�1��G�o�&�����C%��h�w��u�y�`K�pn��y��h�����"wC�n߂�N�\}xx1�̈́�k��� ?#��b���L�z���Qv�/��I�i����v���0��BN�F�%�2����Ą@X�4e���˔%��s݀Eto��*��hcT|�x�T�c�>��C,AJ\
�$��=8BgBBj�D�tp{wh�����������_0v[҅�O�xv{1Qi�n>�w%�I��">�uZw�d~��M`H��U X��!es�k�T�a���y'���_zSrI��Q�8_���F��#�
��"R���md[SuH��f�����@��yW!�TH�S~�5���A��Y�$���}��0��9G1���� �EG�eIoc��0o����2�3 �	T��h�*gQ�E�U�x�H-l�nz�ԇϚ�!�F�f`l�R}1��>����
�1tnC�>�я(�b.A��rз��PO����F+�|���ЧXuD�X�ox.4�&��	�������z��֞�$�&�#E����*��z��FG�6�J��R�>󼢆m��c���-k ��[�j��[��d�@�|%��W�߱akw�L�Z��Қ
ĕ�iWUZ�o��	�Jd�����I��7$D��Lp�c/A���F��l�INpc��Wև�u�Iq�a�=._����uh6��1J�Ss6��8�:�����
�t�aaܫbls��7㑝��N�
�,��n������	Q��,�V�P@�6rv�[t�I���H�ĭC�H��]=���'듃��ʩ�U�?�	6�(t͘s0�?��� hL�7�Z#&�W�1�\�l���8���2��3C]��5�w���(������r���؛р�F�vc���8�����T��E�t�,M��?A�x��?��R�L����4:�Dftpp��ᭁ�m�q�(Lv" bJ�ңk: �5r|��'`�6��t�kS��9�N^Xf�y��ѮI�3������O\���/ �fB��%��k԰�(��,�� �=�Mz��B<�#�tNj���M2�����ٰd�?�@]�~i���y�Y3m(H4GZ3��.����~v���q�2
d���p���Z���לa��o�M�-�^��'���*���Z1�PY�n���JsI�4,.��f1fa��Ɣ+ƪ�$���n�|��B�7$��C9�q&�r�2�UI�Ҭ�V�ov��1 ^�Z$�Ї`l�m,L�0�gJ��Ҵ���6-*�ab{�oo*�)^3�t0�*�7���p�w/MQT���O �X��b��&ժu?X���������=�q��w󉺾2D.Z����y����Ep����܃�+rO�r�PbԨhBw����l��}�E�M|
��?�\,;��~$X���1���olD-�Xj<�/T�*���i�������e��o�7�ԛ���O��z��{;i���kzԶhnD��q�H���0��	Y�N����H�)���c�t���p7T����gF��=�?�Φ��AA����+�k������G��/�b
�q5}A���$����)��9�xf	/Y���)#��{��-:tg�Q���(�6o��΄Ü�?o0j֙�Aګh��"M ���OoAy2Y�+г���񔙶���d^ .�K%��u��w�3_t�>�������$l����M��i���E������V�����ը$E���0�7�*=��(���A��z������=*U���/FJ4���֜!Mx��:��"�X���������E �����Q���nj<�6nd�U|g8�yw�W{Pgf+�R�,�_d=#��=��°� �_�j�'D��8�����
½ꥎ��wﬗ~p��N�E{��s��I��@�y�prs���ZN�?���^���z�X�Q��!ɛ;�Δ����Y2��}E;p�8ȃ�4e�7��E?#�Q}!��m�h
M�?����2��!�-B���ky��$/^�2
Z��6{��w�qP�Z�4z�;h��ϗBm�%����Ձ<y!kA��R8TP�8e���TG�A��,��l2Q���!���K�������+��FO�I��o��}�r>w�[4��?%�'��� RpN����nT,P;~��N���֋��9I�2&*�?�|2���	�\j�9�B�$�]��C�S�w��MDKD��]�o��1��oKd�[K���q.���t�r�(��r"D��x���Ѫ�]'����M��$i×�J;1�&�'$�j�our�q)&�V�5>yc��z�syhe��s���W�$�*���ń��,�)O�cMM �鱖���wT�
�z�s��h��+(�R����<�0G�T<�\-�{�WI��	��㼯[�l�f��j��g��K��1Ͷ@\�o���$��۾}W�C�b�CL��-*[X0�^2a�f������J��5J;��.p>�*��_f~x"EKWP��6qS��J+h=-i,�5���Ò�T$���փ��!��O}�97;7�[U�SAfZ�v��^��r>��{&�S;�%</�@��(:�R*��>�)2M��L�mq!r���͒R2��Le���oP*�h:����4"L/yD(�TH�I���H?�;ϱv���{��	�*�e1�H Y}����`�:�'�	M�q�I!�v�F�)�}P�M���k7�N��?3���B��T�s�<c�� ���mL��7x(��i��������ޘ��%�����ͼ����~O�T��5h��-eA	M�O��@�:�x�ӌ��cĎ��]�.������TeP����ӱ�'��]ta��.d+8Ƶ��gv��r�)��o��U
ߋ�։zY�z�=�����<�ݞcȭ�2���~�0y���O���:�u����vD��o��������� �ߤ�	W��!�Z#V'D�Hvٝ�"/�v-j�:M�J�SK(�9;���[�L{͗��`�m՛�S���=���z�/���X�Q�QV���aM�v�Z�����MMw2��`����80�����pX���J(��)����Ä��v<,S��T�O�D���MJ������Ĳ��aq���5(v.�֕jId�ʹk6��LB/ �S/I�0�k������w��2f|>m;��Ʌ�ʶ�<IO��&�pk���ݚ�~�픎Dz3K��jϿv���d{$͕�+B5�����!����IP��H���gv�/�|AN)�͉�5Y��ߠ�j
"�@�<j
0b !��c��P����V�{�������[�X+]&��R��C�kw��Z�UX�,=i^�-���*c�kr/�챲:��J^�f5�^oD�h��oB,���L{I�9�@q�\�\f���-���f5��{��=D#�yԐ�h��-B��ka�pU� a��ET��w�c]Kݏ�:M+U�^Y��N�(�*.$Ie����B˨�}* �"�r�>�Ơ�S��$��b6,�bmH����Y���}!%������x
���(��re'�:u�ENVs�}���VK�Hn�\_�J�?�ZE� a-W���g�H_|��tGJ��;��"wg2�:_K3OR�ve�hPr���4���c�f'�~��V���˨��fֻW�.��Q�!:��Re;[�B�@�_��V��‭a�2�cAK��G����c���ʨ�/?�G�"c3���q���l��a?o��?y���,� 9kX�1�m�����3�g
i��ez�#�*�B��ɚ�l�C�.��[�?!8�g�/�d�i��}�4���b<,s\�e_�ur�`UÜ�$ߣ�M���=��R۵�V��f������W��d�jaON�5�/H��˞^輝��L$ʯ�
Z�aʎ��Cz< DQ���0'u�M�#���"U�r̰-9�4e
��A罸ʨ/�Q� `��$�54�)r����!-�;DN_�����#3cv���I��ͥ����SM�<:C>ܞ�i@3�Vzzj�м�'(�K�F ��aM��'ϟ��H�:�C�SL�~���%/R3�o��[��R��Gߪ���aa�zUd݁$:P�~:ߺ��kc�K����Xh��#�6���� "��u=xY'fm�u�MkIޗl0�|D�6R���QB�����wr-�I�4䖜�������%�3�C��0̴0��&j*�=���G�C�����F�S䯙�+�۽�B�"V��_nm�_gBd��@��@~���&8��� l8/�:I�]Ki�6p9�B�E���C���O�.D%<W7���Ϣí�sO����b���e�8T�g�Jv�bs�S��ž夥�m�±A�	���`�e3q��x�C �HDiyq�@v�%.�������K�h��+ؽg���v(�g���%tz��lZ��t�!��.l�
ڪ19}�;�09H8�dS�h	LQ�YC����iU����D�����w(.S��%y�ض=c��Cq����d��IR�����e�y��3T��H�mhH2���r?in�C�k��N�DN�ޞxB:����P����{˹V�K����N����"�H>��D�	*$���}�\r;�or��"�=�q�Ԧ=j���x�5i��n%�n�.&K?��T�Kӱ�Ы���n4���O�8�~x���/y�L��������]3����)�&2\=Ց?6�q�����6mgŪ­UI�a�52S
��d=�H��(!� � �|J\�bz\��Ȱn�E�+�乚G8�O4�s���(W�]xeU�^m7�.�M�t�Y=8b��=��d���x�T�6a����S���D#1�m��
�t�k�����l�_@dO]�:�s�jrԦ��ީ���"��ߚ�p�1C����nQ����}v�-����Ye�䵬������jO�4��m����u��H��i�m�̱گ��r���.E�5�Z�!�.;�6q�[�׶�%UE�O\��2�S&�iSuF�<u�3tE��s=g���iV!t�,A:P��/3Tb�U�L�36�roN�<<n�~%�Z�W�:��z��$wyz�����b�>�A�9��GU�|Y�Ywq�p��Xx�?�6�~�}��5IF�y4F�cw#L����:���bb�1P��K"�8[���������%�[8�	�-۲�����Ԫ!!�:�� ������6f�6r)P55�bo��0�̛�ȴ&cH�(m�J�Q1��~����s�:2�q�|T���+1�2�2b/~k�F��K,�&�uYú�:�&�����K����/Hi>>6��j�+)��gЌP�=��P}�=У���+�yC��@��"�̷��(j�{�KL�=�]b<����5MN�L7�{���yf���J6m����,��(��"�PxU�	����mg�U�$�>1��v��2=���h��<Ċ���>����g�d��a �h��	W�/�5�E�і+/(��/�n�x=R�R�ެ�����>�g/��1����<zϲ$�'���X�ݴ��!.����i5�����ϰ�{��x�C���$����|V�8w%�s�
�������ؔ��N���y lѭ��W?c����N4� ��s�>}�׎��`0�f�p��W�j#����c�߭�T�%��<�P���y;���;X���I� ض��ǘ}�@�4����P�U(j�%�"9���sD�9`J[z�s����th�!�A��?�_�T���#B8���yO�����{��t��1N���D?�c�H��#�R��w!_�$4����Q�������Hi4���Df������N'�Ǵ�|��_+B�h<e&giU�|�eg���D^8���#�#=���)� �%B8�֖�c�3Pфv�T{����n���pyr��M���W"x�쐔5���-�<P�%�ܕ1����f�S�v�M��=��|e��e�c{�N �TH�e*Ie]�9gԠ��>Xj���/��V�,2jK�I�y5`�Q�;I���	�g�oү�5F�v����BfH}8X�������
����P��p���r)���	S��\��F���̓:�����Q�sΦV����WA`b'�����3�A��G��,���r��c�;,�q�۸��*Ž�)�s�H�"��ew��Hҥ�R���L���Ϳ7x�η{ey�z_S=;�Hx���th�EJ&Ñ�(�0�Wz`��⭄~�U�D���j�N"����Rm���o�����po�Oku�O�S�I��ݪ��p�v�T�<���D� s���l;�8�ߘ����L���%$#?x�#��M*��14��|F�4ֽ}��
���OCx��f;w���P�I�ܾ(G��\l�gK�����uR�}������K�I���Jo�β��h��E�!�!���.P.b��N����è@�pj��ݏ�:�N/���g�C�@&e�k��X�:�.Q�d�~{j����q�?v%?K4��>���?� �V�f�h�9�q{��b\Z&j@�&�q�s�%B_��W,dh�4#"�u�2V����8�q��J7�'��9y~|&<��(!궾�%��%Rv����E�(�>y�
ߒua'�!��{a���!O_�DB���B��L��b#e�V��1{��S�������ƺ�xv]��}qr�#���^��$�?p�0T��pEk*�߶m�{�m�	u���K��h�Y4��*���3"I6�K$�_t��j�`}Ӣ������&t�-��,�p&�K�1YH�bbK�y��D�L�W�- *�$�G㫲>���E�'�h�)M �1�!6c��O:S,�5x ���Yg/٩o�IpN������F>��_�{�ih����ګr�DS�����I�fX�dx(�m�$k:�7�[���ԇ�{J��Љ�u��̕����e��y�a8�a%�����u��U�F�xR���K{�W���>�+��<B�h�Me��P�|���༾b��Ʃ���ʪ샖��	~p��k*(�7�o��.�/����]��/?�ӟ�:<�S"c�wÑ��=���4گ��i�=����*g�D�	�(��aп�a�>���ȹI�٠ܖ��N`�@��*y��Ԇ�0�^]>jdI����u��:��6��Z��J�hG}�g��nY�r.4�6�ᴛ��֚?٧�>_�$�c��,eA0�Zw���FO|��Hq�t�L8�=eE�F>MYe��z�<%o�a��;��"N��?v�/���Q¼4V��Ե� 38f@�d�DOA�+v���0"���Z_s�f+ߓ�z��Usޟ�R����ȇ4Bx=�p����+*�)�K�IW��A��|X�O����S9��k�p�v �/�ԙϩ���e#4Wi����
���NQ|9���|%|�J���/�m�ǎK��6bOCW�X�_Q��^��u*���<�sRY�,K���˚v9�g3��������Ҏ���ݦ��R���]9���:�]���Z���/i/H(����s��PQ��h-��@qM����ҍ;©��7��~��l�&ݘ��UiX�*�Ӊnr|���JG�l�3)Zұ�.�T���*�+�ZrJ����=������y�D�����QR�S�lD�f܇^�Ǯ)8;��=�(,�����z>f@���w=��ϊy�2G��kB@b��lE�LZmV(zfv⍙?V�hy"�M�~���k�?r�����K�KΒ��(�e'�,�Ǎk�%n?�OL�Dq�� -����|���L~��\s��&��w���(_�(�H�&c>_�N��T8�T���Y�Òӓ<%��5�T�ǧ�\ݙ���]Q���Cx/������G�k�9���Gsk^v�|�\�?Y���ƁF�8F/�Q�hH�
,Q���9M�H'��G�->�����~ׇ�Y8ٽ,#2���?��=���u���~\!���T|G�y��� 4�n��&���t�I:m���f�WI�i���jP��jy1}ܬ��!N|�"4ҧ�\�r*���҃��&����+>҃�jL��"E��b�1�!Aʈ蜬}m</�ӧ�q���w�N�i=>���c"t���R���Y=�m�}�E�Ҋ{�U�`�M(�d|���2wiϔ�7����h�V�N{����ԮH�p���z/�ͬB�s`��5�4��ă��8?�� ������]����+H;)��"�!s,�K�����[���e>x��'@��:�.z�p��sC\���C�����o{��yU��dFp"�_������ T��L;�)p��۪g�g*���Q��^�u��C��[,Z�x��zy���q���͋��	Q}�������T�哆J��'�������cpbG��._h���m��9��T��q5�Y8���(s�գ)G���^.QI>{�1������S���(c��ŋAĬ�dbQ�����e`�J����Y*�Ej�)����Ck�ƎT�-��L<��'h �ԩ�u��p��̛�����6G��l�c��ZKVȀ��~̣��QC��h��������+�s�*���gO�uAn��EF�o6�C�A���-Y4�c�JY.���{��[�)�
dh�����z,�����8V|~�f���rٖG,���L�}�9�A�T@=a%k��q�1G��q��"�����ޒ16������	@lx�{���<��4�E��[͑ "Fh���􇰝o�\r�{ʒ��η|+��]�N�H���Z-�A�j+Kqw+B�{�3Z�ϵ�͞�a���8�g������
����	q�K���"��V��L{�=ϋq5���H:��k�_L�@N�c�uԣ=�-�좧D��7qPu��T��ZQ�j���OH��0'�b�$��%
����C��8.ɣ�R⍔d�X�o "�xOo�W�)6�x�Vx�a!�dA]虬�Á��*4_�a�0�"�>���F�V"T{m2�z1�+��υ�D�� ��߭�懍i����D��5��b��AP ).���M������ւ)�gX���W��;�՗5���I�a�#��l�$���ێ�$��¸\��D����v>x5{��qtw��q_��C;�����?�Bq�<ȶ��[�|�����D�o�xlQ�A�DP�H��w�<�an5�yN�N�@�K;6�ɣ�I$��]A�%H/v�m�����mܐ�HW�J����tܖ��U��g�y�^!�W��қA-�#�[f{M�H��F������b��L����'�}�|Ջm���iM"H�b�<��G�
!��z�
&��B�z8}H�4+�E��"m�������i)����x����_g����[3���[����"���l��`�I��_G?�WP�M��BA���@��f��|����))�c�Τ��MF���� �@r[���b�*j�6w��"����s�Y��9���)�|9
<��λF}jD��ud��̐��)�^,J����*���`Rd�A� ._ZP��B�+���;ɚ�H��s���*�!��>_ʯqY_\���5���
����7Yu��sdߎ�IF�"�*�F��Jj���A9��L�؄t@0��ӭYs]@R^Z�U��C�����B��@+��2�#j�4J]���7>/�@E��U�Ag��ʉ)~��Z�>i% ��\�wnub��dZ������$Ù��6��L��������oL��M��QD���V`�H�."M���&�-Rܞ �i)O\s�$�K�[b��s�[WE���I�`;)T�V!t��6��&g�����1�%�H����W��CǨ`KtiE_����S��}�S�TӣA�m����U�~|��M��\0Db��rQd����u"x�Ѹ�{cHן�t<P��o)=��ds�~��_I��"�6<�*r��m!Nۙ��e+�с��A2+*�T�N���y�p⋐'���û��s7��@e|������0�7���'z�%\^6�~�0	mg,�2>�0p��J9��Ǿ:�Ι��ʗp�{@7��n:�y���x���{8>�fq�37	�(�*:����6|5�$5���+�zH�g��&@Q�qi	�7�qR['b+JJ\9:�-`'0"�|��q��:��Y�S+���b��a=�q>U�$L���G������W�!=}�T����[�'�����T��bV�tg[L��J��K�����G�Ն�`ic�I<� ��(����T0��U%���:(�"��q����M'/aȪ�X�Xrf��ꅠ�6Z^b;S�U�gF+�j�)���1�CTV�h
M�:��䞗#�fs_1��<RH�En9؀BR�f'`���T-��=aх^�1W�hϑK0��=	�u��*�gh,͔�n�*���"��k���#G�l�d�x�H�) �@!��Wed��c��5���c���Z�l+f�l�M��X��lJM/�� s��^2/
���j���ho���HY�L�p��DI4B���Kp����i`�ǿ�5�K4g���8�ʔ��7r�~�P�X�9@-Q�{��b8ݖ��uX@�À쓭����gK��������ej������$ɏ~�����Ҹ�1��,rV��Z/w�Q�a-���a�h��,^̲��4���2�R�Qz� �T��k\��kA��kA�dF_Y%Nck3���2���G��^k�W_���{��gx~x��Up�	�䪬$W��Z2&,QYD�1�I�;jm)%�+�O�Qp��n��=������Ob)������U�����1m
�	0��n���P-�OB��T-P���ö2߻��u�ul�]��s��|�~'ƪ��2ܸ�`+*�追U����H����_*T(�{;��;\_�'��f��"Kҍm�#bY�n��-�`��^�T�ˁ˓�7G[���������θ�sWεWe�A�9@9f�$���"�Q(��g�kD݆�ڣ�d�-=�J�>�64�Ds!�0�j��a�z�<U�％�s�0��k����I�㻺���}�r4�I�=��~�E��y>	��@�z��
f� Y��ö�t�Fo?��l��u���+&i��Yj�x���Z[-����טa�L�v;-�|��B"��CQ#�X��MN���uy���z�f�<��Mͳ�1�h#?�s	-p+n$&y�����7nqWK�RC���Y�$^�iQ6T�G�h�
��g:4��]�8*,��ҬO�~�r��ۚJіغV2cD���5��V^�ܴ�`RZ9;
��G��r��iS'w�&�G�6�SC��y��Ij?��\/P��G�|bTݠa�y�6�yV�j�d�!&ǩ�^Y
3��ݵ�?'e�cH�iPz������J|�L,'�AL���F�l�����K��s)��I��6���Ѻ�|���&�[B���tҨ�����0�R�1xf�,'<٢	["���K�n�=l|ǵM��e{VAǠ�ptd�����p ��"x0����S}��l�)�q0@������������舛=y�;�-_�+��#whF�<��Q���M���7t�LɁ���pp,cϿSeB��,˅��@U�ɋL4�ܡD�E��=�����4�(�-0M�V��Z�R�i���r�F�21�eQ�z�l[R��~�H��N��L,n-�����a�J*x&���L�v��P�J���2s.1��!���݇;&*���=����T��C{P�oG��7fv���?Q_A���t�u�t�γ0��}�7鰨*l�;e!����Q��pZ�{O�"�h���Ir]��x.��{?0���� e�vu>a������H?�6�8Ig������K��l5��r��� c�@� -y�-�Xdۏ����<J�\�����#�h�0\�9����{�$�?�x� =���ُ#u�����w�;��J�m0(�c!�t�ʍ qnȉZ��R��J*W%L��F��Y������vh�kv�E�%/��\�Ǿ9�$���o����������A�obð�K�G�(��5���\�o&Z7+s���[��(_�g���5`�4��9Ó���xQJ�x�Z��,�;b���\_�H�y��n)h�DʖxG�
�& BZ�(���C��"�ƪ�,��G�����>m/b|�%��{д�#���߽õ�tY��<yM2�KG��O�ѝ�8�˘+�!�֣r�`�_�t&����8a+�zjO�u8�3]&��-RKR!��i���d�x��^=Ɵ�H��ٌ�z��WZk�I��)F�x5��xt���1c__��MRbC�v]Z|L�}��8y�:��wc��4��I����Y��w�Q�	���^�U\�������r�84K#�HA��)Fʚ]j�p ,��1Y�Y��i�ɔ�x�W~_�0�;�G���ɴ��P��]d|\t4)&0��ᵋg�����
>�|
�g��=�Z�T�=n{���]�t���T�������t-`���~x
aDa,�L����T�<�]�iH�:lM}C����##�&��~;��QEJa��EuF�V���#���L�.޾�`I�E7[����F/,v#u��	�|~NЕ�K)uT����-�A���2�9���v�	�Am |�Jj�ӏK�7�>!��Bi*8� N�sġ�u��.��>����8�,ް9���/�w*F����2��E�1tf� ��J���93߃����֫)u���:4'6���Ĕ��bGdiS����|��n� +mw#����zAܙ́qF��j7N�%��C5��j7>5��:Y%�}9�}�� T<�뛖�&Ro��HO���Ez�K�����ؒ	O��O��cQX|�8W�!�aXyö%�΀�jg���ё�=��sҚE�OxAFΌ &=	��@w�5�NŹ�ty0����:D��\i���!�y���a�W�3"L,��){�y^s��]E�9;%<�1@�B+R��c E��9�� ��p����F�Ll�Ř7���RB@���"��*�9*��wFP���P9Ն=�S����ݠ��x*j�M�<���~Y���rMY�ߤCH~�*�,]�����u8�!,��`��HUI�0.��0L��R�Ԛ�t���G�'5`�{#p�
�6[6�p��v��edDD�9X��(T�-cr�A���ɒ9_���9���8n��ڇ�|=
��S���%i��D��De�k?C5]3.�/����k�/�?'.�v�!)�������s�g*�f��0��J��+���	� ���h��)���^凊�b��C#)7(RME��X��}�Y�B�Q�o\��nh��������-�{>`�8!ыM�@��2�@���������SbظO�:.����__҂G���Z�3cN�� LE��n::�^T�*as!�8E����s'v�{h�L��o�b��1���Wq6D!(��pj8F���۹��.���qKuCUV�n��F����JQ���X���`��_g���#HcY�6�R�Q���#���zo�����m�To��yuJ��t33,��ʔI�\�_g>߂iK��1�'w���m�J/���ؤ;I?/>hm��_R�\�E0A����ȩ{C���^�İ��[�X7�C\�q&g*���Qº���r��ޢ"������=f2{���m����I_êz�X����j*h�=u5M�#�1�ݸR%�DԇUT �ƢN��1YZ�/}��c���/H�",2,g�ѧ��f\����|P�Pǒ1���n���'������]d{���4�M��N�h�	M�>ƾ�-�$�GG	��ޤ�N�j�w�r�n�`�D�߾��l�A�v:]� ҹ��$?a
1���ׁn�N�kN��Um�QgY 20�ec��-�	��#�,L;}S�[~��i^=�S����i�����6cuqp�q��Uy
�3V� $��ɑ� ��-(q��U�ud)�$k��y�a\�m��$*��XR�;�[qy�`��:��B*�F��/�@���|��W+�W�@�|5�칓��c�S)i[[[��tx�.�A������t������le���,t^]��6����0�E0���*@Q���X1FZ�^� �U��K)|1l�~�Q�n.b$ʧ����wMFмb��i���K�C�)�5V����1������g4��[xR��-�L+B��C�m�xM,I���8
��A�J���+�����ZZz�P�� ݪN���^P,�;PE�1)l٤d��	v�s����#3j�i��j_�D7�.3�OL_t�HA�_��&�a;�M;m2(}����\�<w�u�k��@�W	�I�r3�^�9�o���#:�Φ7WZ�:��3�/C�k��L����Ԣ�l>��y�g���yQ�ե(U��޿:]m؜-�@hܜ�G�L�jA�*+U�+��������q�����d/��Ig�:��ۻw��Áf��E��	��'c�k��r��\�.ܘ�1�užk}��2����_V�L���Qj���Ev�;Ι��uky>� v��<��8�V[�y��%�{$�L�{��j�����ӭ/�Zckn	����-�N�@K������+�~��t��ps~�ۘ���!���:M�9��2'J�)����bt��w�&0�����2����_ș�I�L�}�w����pّ`Ln�bu�cJ�z�O��T�1�#�Ƒ:rk=��<{I�5�JC9
�l~Z��Y��萾+T��-��p���G-��N���2�S��(1�t)�P��m��6R|�O2��k��\�3.G�������ӹ<��ѯ'��u\ww�H�r1����Y�P3&���T.�E���{t`�R�\����]��p$����#P�{S_���XaVq;̢n���!9��I����A)u��?h��ǯ\��u�Р�KD,T'�B�r�����f."3z�b�����������M��c�t7��E�v���<�*�yYe�x�@o����y�r>������ F��Je"D�r�0�+��$������j�T��dO�:�̬|��}�cx屇�n���M�y�G�6��bІ&`����� ���k��kL�v��G��qC<{Z_�'EoتADZp��� M�U/�-d��Nn���w.αD�"�y-_��y������t2w��׆eP��rZ�L>̍��:`�}�7V�}Z5!a�/ز���쵸($93IS���@bd��x^�`�;]?�ǣ�+̞��:\���y��d�4M���k�X�x� a@�� qw���A*��u_��@ް��z�ֱgxӵ�[�LHLѮ%l�o��jSLnS��&6�X�S�m�����'zH3<���_�TD(1I�=�o{9��}[�!+Z����7EV�떒|�\�q�>h��tnA�h�?K�+> v�Ϝ���`W����g�]�X��O�-娄��Yf?#�j�6�S�]H��	*��>PI�ŝ'#���b�u@Q�_�.�#|��F����񓟛��C��O�>�b���n`t�,�Y�|n��~"t1���b��s_�>��g<���X�9�N�a�sD�@����祺rr�>yc������l*�K���@/��)p�4���|�eԃ6�T~���]Oɳ�ϤRZg�5��z-�)�5������4���6c�t\�	��w�;9ܼ�=[�����������QA�PAA�|��F�W�<�m��ҿBt���X�tx!/��AM2�.�<q��j�wi�����Rc�����#7]��lYkm�w�\}��oi4�W����mD�YT��D�9�K��璓�H,�N�۶�ה�׀�}��Yy�� mK�%�տ,��D�cg���}�ICO���¾^�c���f�������.�ZF_x��ch�f:d`*d:��f��	��׀-�0����}G<:9<5�^��&�U���)�_�/ש�1*@�a�
�2��}/>M�g��Ҏ-)����g��0z��=���)x��Cs󺗻�n���(���ۉ�_�q->��Ϡ�>�������I�:�]B���ĉd�T��OF��ͷD���y�S��;U9�����8ԥN�����ev�쳒��b��F�-v�F��\�L+9��N���$�f�q�Jú�XR�j�Y���������*mS���9m ������T�4a�u��C�\<�r ����Z�ty��"E1䀭���Z������>�YZt`o�ؽNw	 5~�����雦���8�Ҡ+'ؗ@��?\����춛����P��'}g�]l�r�Ǿ��j�B4�S��G�|0�c���A�N7ә���;yJ%����(��ڬ�175��Le�>�3� �EKC����'��\;x��d��8k���a�00�&����0\�
���g�� u��IV�+���\j0�
�	ώ�4ohtYM���\?d�!�9��HOX[Oԩ�A�Ηh�A�����[ݽ'83&��b�_đ0�ھ\�G� ��Ϥ�w��
�,�n�fM,:f�8�OX�YjrI.$�5�����(� �3sT-�<)����y~��C ��a�?��~3��riQK4k7iA�����\ ����UU~D4�p���M"ԍd��޷x��)J,���-����l��1����{~�#:`:a��}�ѿdtZ�Ҽe����Ty3��ˮ�����т���]��9�3#�l�v��މ��"P����'��wo8�������WU������)�՞���K{����!�6��W֨I�dJ����)���%��`�=�d�=����~���4�U�n������G� �˒,�gi5;� ƕO^3��6ϳ1�_əK���#���FS��к�H�
�݀�F��9B�i#\?o��p�h�wW��iCH �V�����Y��w��Pi�8�56f(#k�c���7>��.̓��l��J��NY�^��i�&����� sFj�s`Nt�\��R�,)B�F���d�s"�g�5b d�p�����f$�=�6hU�0i���� �W�Mq/w��W��3�Q��9����I�I��A6qT�KQ�[���EA��j��t��w���� ���fR�2�>�²)��	���}F��ږ%���I(�+^X�*+���R�Q�;��d�������9N!+$�>�d�˧�ێ�ep�BN�Esm�S�2��p4J�O��^��ZG�v9�!�:a�+�7�F�2<��`i��=�=_��8(�'�.���4��'��$��SM�(C�3�6E�Wn���#T��I�ϳ\otS 0e��9���'JY�`��7��M������G�)��n�f(�oW�umھ+=�lNxY@�2gN���nן�2}����d��I�;=~隷&Jhx���'�&�YQ'��a�ǌ Us5����Z�a�z��m�<�_�����c��{p˴��B%| &ROs���`�S��ü�U·�aFǈ1�ʏ�Y=�t�S�w3�4�J:�1��\������PQ�!v� p"��M������cP��6l�����;`�b�;�5���ts2~���rr^&�q���؛*5��A�C��h�b�4��[��	Z�_pZn��^�Zʣ��S��G����7�v�H��o��O� p�G?H�QK�ܑ�,|=Gn=QW<�d�LV�׭�A����b����q��� �NSU���w��Jo��l*LYwZ��_�欭�3b���N���+D���s�n�2������s�%�-�����(o��U����;�4��^�$������2����ҹ+(�ʩҏY��Y)\;r�-�G������=t�}����>j)+#!�|>e8ysǅ��`��C����K�:�F�Oi�A�S_g�1�x�$��q#�Q[A7!��#6z�bz���>j�{���Q�5���HsЌHdFAk�}$A�W�V�����T�)�$`p�	���Y�m��竭0���cg9_~@о?����GLF�t�.=��HN)�n�另�ذ�3�x�e6�8=�8��E��k7�"o�
��s/e�K�֥�Y>��Wx33����=��N�v=�S��M3�qc�������ѳ![q����S�G�Ň "�ir1'�<���H���� ����i�wj��R�r�:Km>wL���ƌ T�U������[��� �{&z�uH����$�eYJxa�/d����蠆�9���h׽?���Y���eز��D.�5�ݝ�u�Vj�늏8]Pat+S�E�0u8��m���WD�ױ��-�e5R���,aO�3���B}�Sp-�D�<�A$n��֥[d����;�S�IJl�A�r�n�<�t�����-ߗTi� �6�C~D��d���ڱB������[`�5Z�)��Fjfv�@��Y5z<������iJ�שS��\�����%]�6*C�~�[�Ka��j�)�~�g�%�^m:��j�F�Z{sC'T��C�z0���Q�/H+�>1�*m�dm�f�aϥ|� ���AJ��m�<�1`f �,Y�%$/�*Ξ�8����'^�RM��2�|�P���{��h�e��e6���Bi0d�������`�m=��:x6��r;\.���[�\��~��|>Ry��cd���7.u��N=y'T��G��0 ��/���e�$7�<9�5��\
��Y7Ml��V2C[���*;��K��:OB��w| �2��S뇀2��;6�P�9�:{���H�p!��574��%Apnt�$�2Ov<E���ۑ�3 �:?�y��w>_�O@Aѐ�Yn��a{���[C�O��A*,&�
m�M�knC��G�{�n`H���		'mې� �~"���KХ~��ڟ��gt��q]�K�|�aRv(K
������[��nm}���rֲ���ŧ��-�8Ҭ�D�xbCV4|[�8���|��	eI�̾f9�6��]�є7]�L:� �*rT��Gڷ:ct�!�LT��sJXvm���.�؂��5����dr b���	_�֛�A�|�L"֥Yw�Ū�2�#y��UyJ�����)?uϪG�A	�����r��> #���Z�]�l�(��e=�2��s���ȑ�����ܟo�%ȼ!mZצ�sO!���Os(]�Y��c���{.ld���R�vq%FPN������Tb<m!�-B�M�5�0#�� *��
(��,@X�e��Z��"kpH�٩�z��N�їV)$�lCb�,��"%u�gpd�hOb81��#oJ�^�x Z�b�7[��əbo��"-Q�9,%V�c��ޚo|[�#�S4_D�{o1a6���/�@V��`j���^ٰ��*��2��x̡����XLXD�h�@�˰\��f��S��h��NpX�B�Y���%�W��4�ϭ�d�
�-}Ld6��;��f��l,q9��C�EF$u˖�z�oc
 �aa���F-�^��~}[�_p��^W��ٮ�*��)���E(���(�.,����k�X�h��xb����F���E�xs�l��DE ��j��_�Ie�?�̲2�Hߔȇ2 _e9>��1h(���򰫙;Hм^�!9H݌_R'��qJf7�$'����	��J�߄�h��ԟU�U�iԶA��W�UA��x����^�1��s�I�Ey�������a�r:��D���s����H����v��,�[������
b�T�K��oN��J*�ޛe`�3,�@( ʹ�x^ς"��Pq�e<-v{L�|���(y��LOa�|��=F��@�Y����~ꍅ��EW�߲W�$������7K��;3�-Bf�G����i�O��ҏ#�i_i��X���|�%bO;�gtQ�>���la�d��c����۳�a8�U�U]�a��)��y&8�� � ��(�g69��U��Ņ��о1|ی>w�P��"�2�Zx���O����xtP��!D��o�T��;����*��e�<\�/F�9���(�D���Z�[��#��)���61O�Ď���"kkO4�?���	���矝
]�`l�@�i���w�-�^($�͙��t�`ߧ3Kև�C��4��d��<�Q�Nf`��hN����}P
�U��Ov^]��F�ז��������m�a�4�ޭ/Fvf[�Q�b��1�>�����%�|��4]"�����N��z��M�T}@���u����|��f��*�#h�Lm��K�P�)ʪQ��9z1[����W�x�#��5�hS�®��e��C���z�}0,&�������OyC�?9����k�������H�4�gJ�t�u��@���&�IQ�l�Ƴa9���H�����2g(���an�[��X���yE0ME��*TJY�s�t�џTث[ʽ����]�K��[j8=���
�p���([ �l7to#^�b��,������?�u�"E�k?����˵����6&#G��V��ʾ�u9X	����'3 ��#Y8��<��o��0UTR�9L5J�; �Sn�i�+�-����*��V�.ЎdbE�"�	'�4�N�47>�X\D�9�ؿ&����?F���F�T��˔(�Ͽ`��Fy/Jg<C�bu&R`]b�H���dw��������ͻ'K�NE]�ٯܙ��0b;�,Ԯ�<m�j�A��#�_�R_��qt(3O"��H]��:�j1����U�
��g.�(���ШM�T+ʒ�	î���t�9>Jk�E���r��u�.��j2c�?��4j���$g���f��&�}��1$X����f#��ze�����u�ȁ���LX�»��]�;B|��h�ݍِ�}��m����nR=�u�D�Fv��(��`�t��.�y�l˃�(TW���7�94W�4�5���?��>��L���òj�k��n�B�ш�����G�{��*[�s>��]���s�
⦕�@�	�zV�y}���+Q�$ooA�;����MJ%]������ſ�o���u ���k���]o�up|$������!k+�W