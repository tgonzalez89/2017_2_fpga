-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
IyBo0FaLqcJm5QcY5DcJ8zfgdLiggwhM1J4x3Zxxu9LpUMsfWYgudG2labWib4yJ64GdZ4HKDuDb
xz5SSli3NPMyzfRX8FPyVu0aXQZy9en20ILkWiPB6oT9woqCIr19jhkVrdyoYhV25NkrLh8lerca
Zw4kfsCKJK2v/NmRurnpS8K8CHnkEkWm/s3Ma4ts3iKZf4fYfXEWz+8nWLoZcVZVaD/u6JdxauK8
t7TOB157uisarOYw7cpLZ7XUzhig5LkaYmNn4bZ08Y++lMZEFyoZq+k1NPwD1ZySlw8/TgmfpO0f
yKJ3cYzakI0LV5/ajrvnfQprByNiFxQ857hLXQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 24144)
`protect data_block
L9FylX7TpFpYuGFVuAWziRlRNLaD8iSLuqauWNiATgONXEaZK1W2uZ69DYjvY87sDZvKBUXUH3M6
xJ0+wDBCawE0RkMljCwbV137pDotoGz5NMCkCPrbkW4ZOnEz/HonlDzCuEXFSBGoj+O+IyVBZCYP
ABFk3DHUjz/qyxd98mrbWA0Wt4xuQU15BH3UYwXPoIzN/Kkpu9ju/hwzk8TzIzbRqoyApS5de3qS
Rd3/LGsiqgr603or6tlfnKEyDerk5JIrDLgPq424hrUUKug66tfljZ3Oi0IdSI8jXKtvYW2K6rvU
sOa6FxoeJNbbrxp59l2n4KoDzB8POMJGokrEZ+BtRxuz1a5lmLQ6muRP5LOF5N/o7fRcsiEH9lIz
2D25HFy1V7G7YAre79x/eFjQ5moLzp6al7589C74YpS3gM6tlwjWj1qP4n3gsUXOUNIK0Xk0DJ4i
IPxR4md7BtWP3ZcPMfMGJjkjBGKcIXfa0eVrC/cX+NfNiNgp6PkMIY6HC8Rsdo3s7uVEQxLKZQPJ
EPlUCCTi9xizQGbKQRt0jAmq541lmAyiSDdD/41Wie9UaVkrOj2eJs3M2dMRwo7jJUAjsFCVbJE0
Yt+2XLwkQDXWPi/KKl0UZg5GYBHMF/HX2Qpt3X3LtJZbpOC9AdSUM4mxNV/zSbEN1dqxd5QzsuK1
K/tgKPnqHk2dnQjsVqEJ3GUJCrMZRif0lsGKLtfzzq5mCjeYyXuVMrTG2ZJCjyX3b4QCHQ4cXxB+
pZAVp/zlnbfE2iLtq1Qhw3mM8N+rNMqy9QM4N99eyz8paBktcixXxgpCxZrCBLi42rt4K++W3TUZ
rpbwrMVyZ71RxDGv2m2DZlUpWGi3iZfKjWNEZygN/wZzq6XVbjIjgqUnEoc2qlOWbkCQS7EL5CtT
VQ4dI7RlVU420ljcrvnW/PlgDSfbT07rbDb/XX4RkpEp00QgTgEFf4kfpAxKHehL210LKDSbcuQ1
DibxWfqyKaY2YPOpzxL0ptZMfe0AZJ1wy8jZfHiAM7jyNAV56J0wENVfDccgpinR2Pkdh25uF2kz
I/ldc0lwMBEUIkyJlJ4mr5uV9PiobbDRCFLRiOP3GmkgTZ3NIbGiosYjSzKtHW9Nk4ot7At7gAsR
3TW4TRYYbQl4vcIPolU8Oc4mT8yYfwCFP0kE5GjguOjbqnaVxbOIMk4MNOqZPxd2lvtkyPSVKeXC
t3PJ5cEZNkDVEwj/ofUM/1cE2aM27vz5jqTRXUTyXS7TH8OvF+P6yGesLbAZF7bzyczLqZgLxwrp
fXLyNHz1ZSCeEA34gnaIG8zxl+5EBsadpH5G7H6AG7HmcfQst/tofY9PIK6HBa6YaBosPCXHPe4t
tXHZvVDEXgublQCbOiwqMmSN77/SvtJT/WzoIZHjOcT3DjHbNr9OguWOuY9j3l6gjdMMtzCqacog
eAOOROe8er37EoGL2QWmYktX0QZxImSNXB0kTBu2NhSqXtIYjlYpWqIYBN/FH+LhWHWXiEZKvSt8
CA6xHpSpFCOQs8fdSyP0NxnCoPtmAxFKIIx1kGlMxnyXjdu28V6W8gjIA/DQRvRMT5BKQF5g3Z+I
k+//nMYd/IqAsksgMT326Lkw1BHKSQEkvOjGlE3os/ogU8fCucNHtbVK8kGNB0rbyi9gQIe3/5GH
Wikx9ThWwCKHkYSjnDGJ/3us2gwzu7kL6wLDIFiBnJUZukPslKM3WwwXvNv/HSz6qjkPXh0cRH+O
VleRBLtSTftGhZZeFzdbJVUstjr+dTrz0lkKedu1cZz9BG41UxbcfLRjIv2OHaqxAHdElCaAQ6Nq
RxeiRRQotglQWSwoQk++gRX6RgBnwaznEkGh02BVvuddNqAFbrx/CCCqtxxadh6pB1fdn53ai+Rv
YL1t+sVUKkJeMX11sR47L6AJB+XvluAIyFyAvZkJ/1rjzIkFG/WJDOMrKyGOSbHpQ7RmVud7kJQ+
uN1n4HnyF8CxnOc6z+QLdb2uDtUY8rBgI/t8scIAKiis/GC+geLZjWcd7NROVS9K0RplMueNmXY9
g2k6rBVu6BP1q41nxfUU0GKbJBwLvNvAoPuL59XXh/h9l2q5IYYaeMd/PbkrMwvD6kXwp5RIuvFs
bSVXiTyKxrYnTLTY8+Yk0PJ5tBzEzy1Uqhj0FbaqbolsFAM2z2BEPh6yxq6WevafUB4ritn3NrIO
M7zpZUsrYx9k8LryuSyGO23+lYdQdLsMf9xHUOfq7kBeXNQBHzRIZvKkNnwhoqh/WooSG/WiAR3b
3spHRV0oGzOc1ySxqnsj8jUiylcSfzHtjMTZe9FzEJvf/29fvXfC7jFHUhl3BBMw3lZV9T/k4oBU
TgpEW6yTZj2DXdOsviNNa/zwA2M2dgFU4ABaUVunIUULkt9i3KZYXAbsQow0Uai/TbaR++irwsvF
F6rZaU1hU59umrUA3FaVMb93XEz3vu/QBpJJc7cw6bScUgWqt4rzH+dwlaJ0dcvSC8ccQdANkG7G
3dx30uo2wBB3aiFD+yWpU2DwkG9FgQOts50zEWNcNBOsIK336FGyB4Wts4zP727EZdUp6UnZ5DfQ
SBjBAO0b3f8ajBHueN53Bom06v8CHRux3MpyRfvParMfyCiN2CKAo0MaIOqKzmGBRGJ8T8wbLoEH
C9ruVyblD4327mz036y+4cMHZToB+/OtqOnex4LmcLs+xLZRsUr67UFl77/lfidlZkgJEsnu8+6D
FBL+eLYehgFJwZkSU9M20tYK2tfcMbo13Yy1i6fPw6gL3j30ozpsd4qCwefqSFIq5qNDmOKMUKY+
B+XbPieDQASdLow7YPwGX/AXR1/2Fl9/HPFBk8W3pkaNbn0jza6Dp1vUICDYS66nSAD5MViYnaWG
k7JOGVztYWt5FV3Uso91NkojpErhXNepaLLtyBA5/s0oyRG1FWTyw07P51j/z2nOD/0hpJQODByB
GmZtloLJTyfGXKZSJEOKiIjm+jywsVIUxDBpKCMCyDDJjR5ZqhOaRqhsbgxKXQhmUItuhDOjX87d
havcNGpP2YQVrbOJpGBx0duDP+IFqWque70Jrdpzrr++R8lqitv2CQgGA5y1suJyub+JRGzz7W2H
EH5Qn7SJJh8Z3c2WIjf0HmPkwy+pPDzDfQNF3fnEWQw4vYlp+g82xUrmq2vqHuFyaarl0pogD7OT
q5jZA71b+aXHB3KaujprRLsmhKmyho8bF1EQckJ3RMROPbdnGNCmZu1QunbapUk+LjYHmCLi4JK2
ERHZP4sXc4jWqlGBSSFd+4eWmDJ5JKqSza+63GRaXuySUbJA+IIoIYUCnOAMFI+uzrjIHQhAadrI
+qZ2gj15LWFpjQSg2Kuw57Opd1HtVYORJAoPtB3PsQ20QmDeqyVGzXAA/h+ouylspQmcO5GnxXGo
OPpoERRZ9o1Itqy+vLl2Ct3rR1hWvVNDnPo7JgDt9tkA4YIJsD6n4Cy9lJtxOMewojER2Qy4PPt9
d//kY4A4TNg5obe/l1s8AslgIu38gjI2MObDSyXO9rZcFU01qP9OIZBx2MzfGAsjYvZSxPlA+Slx
DiNqHb47BW++JTGK3U+lYEY7mwMDWumCriuKD4tgl4kyTSmpYQPwyl6Bx0Uf7dQSh78oTDFj2WGD
4Cs/XvxDts02Bcy6lYZzhmdKpnYAS1vjTOJEBtwzunVdBXdwCX/JaxG82QV9HDszpt2Xmq3fyA+X
A5GXhnhA/SOqOnK4t5ysQE8bvOMuf9aO7PU/TFuOXXFC1VvzuEpkZVmOu9M5ZNQjOd2eMcXYuaoo
f6NbNy9S9g6MxF4iLIt8uQSmGKCKVRVzRTIISWb/sHHaZ8WxcqMuapTyCkxr47OVwJ8HK9tis2Fu
TxK9i2LKfCFHOfUaLNr0Uh+amoFt32NBC7ukdloj2aXEQWtFvaxHgT1v0fV4xrJpgjYEvem4tog5
0Oef+ZjzXbXThZsfHgW1SoR6MMWBgWSS1PVlo4TPei0H/IN0Rad2HKjuOjHbfEZQzDuxXxI86bES
mxX60sfS7pRTShBXQeZ1XIErfK5TGEbdZowdcy4VX3nLjXaYNOKu08XXw2yDlEQE4f0K4hAq87VI
i+jPaV5K0Rb7ExLoeD2VmMKYi0+Rl1g6258FH26lwmRQh6L8Y9ipEqRoynZvqiX4TWwaE+LMIOOT
lSOYcDokw1H0JEfdkRZyoDWQentoq4xsjTOq85uiS+UTzOzVBuFYy196p8Yy8m0H9/Zu4s0InaKA
XmDr/YzwUUqnM091yMUbjIyP74PdGg74PXR8FE7rLfYJg3yEP2NkIgJEDmjGKEDy2n2mPqyGPDo2
dGTjWjHgeYVV9RYnVrOuTnZJBpXhQ7CLbixgkrPuLkVc1mI9cpBtdWgk2uUOKs7JBEpxxRr2o2F+
e3/0ubSwVWohdPYzBwPdbAUzO2wULr0s6LfqSFqjrlFiXmHV2AL3acOBocW4baCwuhbdnEwGXslN
6+LtX8Wn3g967clHWlpwm68lUMbmJN9EcIcXKGct16XI05NvF/Mzup5X1giESOdbzczLcCZNx+pN
SDTunM3gmrRiN7QqstG6RYNYRtDQWPJV6yx3mKTYigRlrfUbS8UeRmYbErERjOFkZQrFl7Ztwxud
22tMGCmQkF8bsGeJoLSuLbN4GzDUpaOuOTq+Ss1ax11QdYYNMWKlA2NZqpKrJQmsqMnLiYJohhDb
3/rwCdkMrQgbVMQSw4Jv4lJeh0U4T8jrPuilxwJI7Z6LTxMiiAO/aSx1JFjLVwD9NdscxP7XGw4R
QQcu3AQ//0YdxAg6EJWYf9FWbWsOYFmvbycpRBVh7lPH8z6brUCeF/DSCj9BY/KV22heNrOCNuQc
7ww0mzrnNnd7CFQU8MzpZ/rEzK8IZi4+w38b84Bz8F5NXWTQykv5Nx/XiVXqUaMp1RI3OYG7EBsR
sSagOnvz/RsWsjV5gjKI2xuZrEAkuh1zrOjk1rMBlTLkomxM+KNXW0pK/KibaSJu8v94Qt3W7cc6
5+fGe/2V9cIUFb+yc+vSA0ibDGjYJSlJb6QDLS5gGnZWy61GfgH0OLl4KldV6qSplSjWv6d5tiYW
uVa14ekTQqX6k8jXAx7mOX1bDvhRVFsgzq8M3lA3CqwDXs0O38pPZ3e6skWhKx904MwQD7r+SzeI
JMR349CCRDswZdZxsEMk/i84Uky4IzFNkNCbCd3b6iOf8GVrJP8GNcpQ9pRpSZ7z8EuOEUYNPjKn
5hL7k6tIyfdrGxOxCgftvjVYR6sxbiG1tU1ai/ybWY1FWeV29rrwJB2yilJsLlOEBCczZCnj1aD+
Tdjup/RoDKICUmcTbNzWMrXHpJ3ZcKKt6E/oO6rBGUBOZvUISv3U5fIQ7dWrjs3pyUYJWEyiVLu4
HrioMjkKe5KS3efdHahMvepHyk2Rs/qaS/ArrPA6SGu19xXa4OS7nXIUKj3rm/j2ecREuyp8Z/cE
U/gQ6HjE5YXwlhM/Y1+/NJvRmYXH5C01DwXZvWGrblGUjAW7CeTGc8O0McDqWJPYfx2Fxw6KPu8s
ZW0hptG2rutI0WV7dBW+4M4TPRBC89OED0B4gHqbW1kafJd7tfaFaXi4dpQkQx9yS/WQjJzTSRVl
rMUnPYCgC4BVc2M7Wz5Ur3X8VRg2lIEcs37hNwQo4Ow8g4QWh6IGt07jLrNSucv5WDTzSBz2/BPw
hr8+go3EErKv5m4OmX/w5jblGnJkHNUVVDd63TOw6kFhvA732Bh9Xxywj2roSJSwmxLLzssS1u7u
gWxfso0zo2kTgPHrvJ7HGCgLgiwvHLFGPAKZOMHYty9EsO/086k3rUNEHBXO1GnUuW1FRUur4XNc
8N9+9akY17hKqivHTDn5VR3gT+MOB/kHA6RlntGJ++dwNODLL6zT8ki8jowkTC7IQuW+90f/FD/Q
f1vZ7BrBlylWpwL/0vmCjnPOBoKmwYJ++0FfLbNNXfcnlpxKaP6+9FDd5DOOKW8NiNKBuZSIYZKB
hPr3BRXGZOb6NNOjINpYNj8t9SFJn6np6ifSCs1tt0RmJ78U303VXveYbCse+6QDZpzcn9vRaYYN
C2f+G13cE8zpqoUuhHDBgxy0cTJPwDJU6TaeX56r7C9rFUMKMEIfJaUwtCegJ+k6XBngC3TbLDu9
0nYpR/FLubyP33N5tTsESi9W4GPQBTMR739TImAey49Idl/eeus2GltdNflzqND0ZKKM7ku1+ISo
nyYpl98T3+7ZBMiH3YYhTqesoflNr8JTsDtFkhoSXiRRkPWnPKacnb3boHAj19h18fcuZKGtrofy
4z+uS3h6ogGuVJbhztqwPR3sezyDJtBgilZCLOfsCSO3wtS+IBXHKb/2DsR3oJ29pODeJ4QbiXyx
qv5iSLdSp+sEJDQh/ibTrfdTwH9YlPwAeKavK9G6yo/jRNH+pGY3dqxP2nae44appf/8P/u/d28V
JQVugKJTdKoPg/fPezJmw30JyhLp0Mt19dvf3hgffjV5jb3f0oqcs8NGuRTMWY7QNX/NIBlgyYlu
FwG0CMRoCiOlw0GBCpBSWLynYuXV7rhnJV6zkBWl43Gnr2197tAEWWR+A2tHFL56KpqDlRFOc9HD
gO7Q6GHMxBL08NR5AxdcHpLShBF8upW4kCrBkx0L9wz5s0DXN2iudaGkDOmvCc+AWztEHQJ3N4ik
ObU3+5j+meglDWUSwyh8WDy9iPwEebemHr+wizAPEm0IH0Oxd4h6T/i+NXdS9vFGhd6t6fpbYQ6/
bHYQPywb1eBb2njEoeS7vSkndxRyFrpbMQglsDRLSM2L7vyjVeY7CpLE2J40uakZnCPib3+YkIx4
eq9YSiEbCCt51bPf/vFs094CxTlkKryW4uzgkUsYNkQK/WIKMK9oz/4HFO5/wAs3V3lfpZRpW0iQ
r+KaokXZhIL+XvPrIOoQy/QGdes6piSO39cT//8Z+GvV8CeZjC5rIELJ5LwoxPp+ZDWnR0z1p+EY
4N3Aefk5QoC4lZ7du3Rs24H/uB5BfpwgUFS95NOxqwCT5h8sUsRwUAcEtXjSsoYNZQzqGjhTQOKf
FioQWs9XYNzQbAKOo8fnX5emAIeTAMR37bW/wibu3MHCoW89187wWm+rkIHtoK0O0E2l2RHytifF
jY91X0cgMywCcvjunWFEJBLwGT6lm3PMxCUlMulTtkzaheUrNM1u48PbLBr0hpwpO7cuKIc0J4Qp
boQYYMjJWsMqCDcC31Ag2VeHh5vC5kuFzcNAR1XmvgRh6jUCkzMVZ7YOQmnuXCINOXJjBstgXtuv
RGjt5qRKbEJY3vGuVo4apsnJw2iGC8q3eQLkVI3bupZahf7FpOPfvIiYQieIIXdrDmnR+mJwcAwr
ERoS4KynFY6jYSUvkSQLlM0n0Y6dDjh8ruodLChlDaDpUqVctP8OT82wD8mVHEk5ATmnoOd2V7tr
FUc7Ku9+dXLVspdQZU1gA3OwytsTIfJB+kRZoe2YwfThwnDf9fo9MEjG4e9bKyNVgKgwoKJ8Epmy
E5P5OfCNF46/xPK5fjIJfEXl0PnwispYJXyaKY1p2wplw1qneSf2Hi3rL3K4GwRvCSdE5r0LVmQ1
wUQMzbAybq1hEY+M4IdKN89Ap6KbOVSStFUf15mhaXZuHEb/E0Z0RUQLNGOvcjFpEdBxa7qDq/ma
cTgjDPUjqy+vxQwsbemi7MGJlZeKcY4yCHsHfbw5/Rz9WgOCmRV09AtN0y9DNxL4dYZaRMJf/sC5
m/HPLx3oETSaEbhRLycwr7O21KqkkMe/1H+nB6VR9LhxlXkJxXXNhT3opbwBJZi3YfxLVu/OY6PT
EwIcbUJCxGp7gzoKeEnVJo/kjDp1/8mAsZnahPLDXP4OwSucNEoO12f51XLtrGDRFhOmnq4F/bEo
EihF1QQ5RVm1aRzHkuZ0v4rc4+1hMKw3fU/UkHhod4q85UwwOSCIpJQ6sZoJ7CxceBRP+yvGpeaY
lzkLLWNZYyTu7Y2cR/l1JqwRKBkQvL5rspi6HjCT3VpcJm3cSRZGYhAxADaQ0n+iA2TGYd/LOO8l
QulqxzyJLOAqOlB7kftJcK9UgA7zpsSzn8kxSYhTqIz7AQXzW5hMgzIue0/SKr208f88PqmZz78Y
E7ptlKIsZLFJs+kSGoxa+DXzpjs0SZ0hHYQOidJCGTZkM50GtH6BkdR8hgv0Dl2TJsiiBir5ovHW
4sjDJbVkMz/hu2v7xywEXJc4NbzLPltTsiYTgo7PWbwGr9cUVV37whqr+NdSK67rVncLUT5Vc5dX
3CL+pQ5uV1S80RyC8pYRqKZCmFeZKHYhNj+BuCxGn1zxRAHfuLlo8dwaven3u0fwJWXAjDdBngLm
wzXGVEfp3gYdKuE05IYzPeP1nxygmlTUXRHTHYklGCkG9ILhx2pc5yIhtKd1ZhHJ37RZ1rkme5hA
K0J8mrcdmhKedowhFlBSZkLrUyGHwAFRpZJnFPAjZPxt8Woj/nrFPm7VvQyikc7tiR2chSVArAIZ
xmXeco9XzZC0V4WrXvpC5Ds2cnl5i3Hy27RqwPHhRFUrSxIhj87Rr/U8FsKkfqq8meCVb+7dntGI
q7Q6+vJyZ4lWgqyeBju9HOQ6C0/pYPbKBlSTzklRxPOqYsxcWdU26EqXOt0NPXlLb5lLpICvP2n+
1ku2TVLRwnxl3YPsRrij7cdiS77Av53HANVe54BDRvq43pYtuBEQdl7P+DHITTISSr6fsc6R7U1J
iSrHWF0i8RLISvOAmpd8o6ChdvX9En32PXf9l/ZkTp8Tlaw675aNEOQJxjdMm8uHAdXlfDyYBQCW
r56l9VHgK6W5EMdLwC4uSV9EU0ZU+18x4c3JZQWORACs/1M+QuKE2mFfpWXHlvtD0eMyNCerPCAL
g+IbIJ/bELTV7OK5uCFn21il1sXIOBl9+7VwCsiAXi0CRzz3TQGCJJdNOp/91D63qqeJDnlpRzfx
j/COoOCGC2IgmlyeGoV8k9AkMLd/obyPsMNDOmPoqxtlpEQWKV6F1ZOYH4PVxImxDVReCEa2MR9R
7Ywy2gqZGpzuCmLs7xvYBn13LvFKnCHYS0etpc5+tK50KRzy6dVl1wfhwwHmvsXrzTBGPRFFbVU4
FVqlU0rNvQrLO8f4ODqD/WbxB5nRXB82iUgq/Nc9L75F3c0zD5oZ+r8HIhTbzihRxTOHPRTvF6r1
kgXRWm23MTbjWZ38oDXm36gtZJeWSyj4Wt1sq+cxTHr6nxbsFcUAAVNvMB4CUoMRWy7jJWvQFsqe
TyG77lUcj+vpPzqL4rvzZRTmo6XHcRrRUGqoJx/xMLTMJl72e+d1ooysxuN3HtW6mDH8oYCDmNgW
zW4MIcpxRncZW8oY/Q+R8MZ0MMasRl4eNwR34L5T3cY04+RcrwCYO2H0wnTcxiCe3lPSNKGnKVX4
AC86oWOjHBSWUgy1NXMr3gj9ao+0Axifte3Mq2kH+ud7LDZHcV8W4yeIrHgr61qFttQw5JheAZnX
V+/s+3Fw9NBwPLXqDYPFGgisRjljJb5c6ApBCgoJ6p5MY7CiyqEtd4RzwBLU7IZa3pYqbe9cGQzy
crVRlv7QMcgnX7ctiwiUWjkUIhOsZUHnjhK2xMtiI39lO3ONUlJ0jFdbVPNy4d4XyIpBp0ZCLJaC
GfUWeY4IfM7cEgIJpOI/ZSe1Sk+dDHIU4wIMi3bzQMd2HJSakHy8udUjq766iRwjmRCj28hgl7QT
IoQhepcljTWGjmZKeaqFiJV4I2vVH7TEz08X8FOchnvsEW9lfmkX5a15T624Ar5naMGghur3cNbT
q2CICIgT0wq5jk+RxGVe4vkf6iL0/EXWYAiEGql1uHZYDeVEGb6CkLVmSe5lIn/kAkbQ3sQUt17e
PnkylR/DnYMVtGnpahkhodKsWvvxnLqcT//MPJS1lqtS/JggdKqu1RmE5RI3pmGol9jvXwQZ8Mfp
nSKTqtfHBMFSl26R6CrC2YUuXwPg3GR8j3Q2UwLjyF2dPx6Cfae9nEslyGkNaSIgo/w76mhBLtdW
4mrCr7u4kADPlDwSt1IqSGpTksPAwSaj7uTGc1bIqQFvAfVpBKH9WQJ8lXwZQtfur+N0w95VH3Hy
EQ2+J6eXaByWrDUXj9POovaaTap71GrbOyhyO4wfVO3kZLUrlranzrUcJMRklSWevCEeULDj/NIB
aI9BCapBI0dvRDFKTBlBaVw8D6rMWDBpJHD34iKTvaireb742MlAlOaXPRqdGlbthFWnl/nvr1vu
ZBvNkLM3uDobm+Jw0FKtcq0ZMHRxeYt+Q0ll7qiwNsZ3fxSp6h9VFzrh7DeBIc5vfwP/AHZnGazg
kvu2V34dRRBVAGFHVp/iy2S6YuAoBLdWXn8Uy10+AfraIGQA/6Q+KV8b7wYX9OQ0QQ7qJ1tegArm
zSMgg3nj9Nek9LnPVaY5aKD8jVkrN+mqxoFzeYuEiI3Cp41p6Gf0pM88ZrdpXxb5Aq+usd+GVAVO
caLPbqur0oSwJoTUE5lpS9aMR0f/SzLMAFlpEE721xHL0UHeVHb619pqZHF1EDfjqCHnyldEA/wq
SEE9aIP4sHpzeGtVFIrKClpQZgvDoPKg2noDxV5TE0zG4CDfgitA6wQffGyB2GcLD++OLyeuVwvm
acgKY3mk0tcXD1eFVfeN5L8yfzzBXTfDdcXei3xHWwHBni1z6bDbUcD9iEvyGC06dz2EpCw+N+7Z
DjSreGuBiCN8mzFuxYzdY8TWv5J0swriXpLYpLh+9Esoo+A0lmzqJaiW7SzqyySf23zRgvYLIKsU
ahmAC+4byEOKXi+5fLDSn0Q+awdANk2gnCaO1mu6l0ujNrsY4hNZewWPemUNZVZIMilBTB48nKrt
v564Z/Mn4bsoPV9zWs66gFhCObqeuPnEw8DxmtqGlHI0/5HFa7tmj157N4Ujqb9pazdhR+FulKux
MYc3VUDjGRkkrbPVnMiLKHBPM9mKfGWvvl1BSsW41KFX4diFAYXtnjlHGHlXczs51IJm4F+B2wRO
lTO13WJafdZk4mR2Pn2JK5Ox5SFlgqf7YBhT8D9eAMd1MbxQBkbCyLx/5cV5W1irRnuJ199nhq/r
UQgTLn58NhuVrCrhV2UNkBzzwSbgy+0T9vAazwLdee2g88aKDPN6RbJjI68Fn/xRP2PPuQ+YPHn1
mNHpZRsYkYXqyAQCWg1nf6VKKVluombjqRLIkeANzbYysGspII4NQ8UcFihYdGHl/n3mni7Wg+GW
FfH4KOXQUc991b0g/Gacx6h+k7kpVU3U1vusrjWxK7wSO+soLtu+/tbkMgZyn2ISdVg+7DsdHq/W
rjtBl0yS4u+STL+dsiokKh/i0w77tAuCSVxmKETqC8n4svE9mVicSWt8vqIlLcw9btVT0sM3I7wO
LGMlrQto4bg0xjBaTkrzt8IeGrckBPMiaIrv2NWsLGDFzU2f+iJ8bAZQl3F13SRCOXjnbivN0Dtg
EUIOp3MO+xHF6pmzvvqNPMHHqcq4Q9Bsr932aWxE//1VB+uXqv/JZnekOLi5XbVADzTInG76ZGdI
f7c/OV4iq8OlXHTvl1iC7F4S9RVmxINRkylq1V3ZpVDCrq2XCvaKid9AlAK8m9mTQCLo3iXzM69u
KEWCwZtq3BtB3sWRaB7AeuacQ16obLZpQXu4frjVUzw6kJy7JJNjJYpy5kCUMJQJdORXnWOOLQ6h
Gbn+Qd/h1etEAzv9PFYP8jDXj7cqbDJeItwunlg5ao9Gd1zxYIcJXnncYneS36VLfl+/EAV9pNVC
M24R/qUvozGnEJqd0TyirA10SG4CnN/kSJ7j5o5Fd5kfbT8IMw/WDmg/uBwSO86Lrrs6lu6jBxDE
ALFS4SvZKyAJGM7DjTPWbJYeJvCXunUcR62YSAZ5+PJfGdVIFwWd+iJ2zxaNT4JfuVa46GYkZGE3
7dsib0KANR/SaJYfQhyZAu9XgRt9/b7IrWSyGIyVHdu8aWD8jAJwow8K64oMk/E37zI77DWs6qwV
a+LTzpSQTP4E+d8jfcJqJiiMjfe8yC5jfZOJ7Oso7rBCH8jCon52shLr3GZqUYUqvarRngI24I4j
DC9UMYEiCDs4tYaTznHt0kIBxfDGKM5BQomyn0Xc++BHS7PDbJsTi1CcHxc82qD42WTxF0E1ae91
cOQA9wAwJatiqo/vas/YFgnNTRg0gp5ugLFFLOLtnIrfDaCM3rh3zihuaA+rUxmWJRvCPvC/RPaS
0WcNl+hHW5JaU73FJMTGrjB8lhp2WtPqwXGbU8dnXIVJ8UjNgbOZGNLl+u8DXYBwzSRzEcIWHi8o
g1zYqNI+iiIdq9gnO9RQ+yH67AKrbswY7TnuV+MRE36FIWHAJpwErlXvfqbtP5RnvGeRtmx/QTQx
vIwbZjvdg9FtMfxxK+WmYMm0pzwvguulU9pCLqj4SUgAn+iL23hPFrzA8ntK94gEvH2IU4FDNGlf
W52X0wD8CKXPGpSryPqwEkfBwwy4Hxc7+bJy8sWmSYlBOG5zt0MqV68atg9Sot8Tz92UrM704vOc
a1fgKZRkf8n+uD1NEr9GRSwMEQId48Jz5ycqSBilFVhTGmYAJ/y71KRnMJWeKV1vpzyfcH0ZXsYI
wpSHRYAYftw2L3afC0PBugDfCMo3oUL2P2rBv7n7NIvKbgw2Y/vdU0VtUIzsPcH1rxRUq+L8VijV
z/tWJzUW10GZCTu2EVPYXaRbHVAW1bCehnnKfszwob+1YtoHsfYIFykrzVwMNICGmGpYigmfRONf
fGae5z4cG5I71faY+61Y666TRVD4/zAp22tzYNJoYsJB56QLurhilaKV5NGk839JMH2ecfEPRhTP
p6MN2RruN2/hWMqUiDF/SBK6k73ZwJlQ8AxKlB9fu9KZwI6YqJ3vbTySzHlzNJT197nEod4L8wfS
FGX8fNTgvtl3kwbLCbSwi49vBxboV8vPfAQF4BR7TwKck1nPXfhwXJ+7HU2oIfNDu4zFhIhUFWtJ
cTnDqkLCuqZibFk4+hf8ipQ/Z5foQ7a20HSB2nd1C73mGOBazKOMUbv9w0A3XJe7xZCtSG3Quzu+
PA8t6NuFgUwTbMHjTvNolW4qL5LK4zjAAB2KYDd3g7JFqWv0H6dTomUBKe3zk33X/81dudOX2MNl
t3YlwUsYwWBgUs8x1X9Z9PlZhag0Xr4CeFJhDFBTElB1OOwnemhu2FxrDT2sSJEOKNXZeBai/bwd
KGHJGh6sswRfJ8WWq6MOwXgAXSyIw7cp2EkW02opS3xpv85CBIoitmgvYDEyn9IcJsfoR3ww2eA6
KT8G14/FUmBPYo5oAhTiO7u/OIiGp7wO2tgYCAzpKZ+jKzZ5On83QC7Htpvbk6cB4Iww7ZD34QcW
IjcBhRgo6txJ6fg6QcwJySUZM51T2OcH8bt1UdoDFrI43/nojwdwI+Q7hJaNjsi8C3CxokJ/TMQP
0fkr4RrcVmSCn/7WK53e7BLt+90cGIKY+VcIGhgNVXyIya0fvucf+Mq1LhnmPDFepfPy1YDzcKNl
Ydj9/wHKazMTDGZCOu3q60zGvOF9di3zSVlFrmhyabqM5VK8b8FNwU4+FpN9iuQu0XfG9/16kKyI
CptQ8ltFYOYBQF5HW2w75bNirb8ZFKoU20u+KLReMoQRdv9/JkJVeK2c63CzzGfj0u6jHraPGtUa
NdOtiRqYdVRjPwEcMkS7NeftIaS7F+QIn5eVu++zrua0Cl3hZa0Dw9MuQ19oeZmE7gTqg4NeaQbc
tyuGOg9Zo6Kz34tbCY13jQfpP7cWo/m9zCpSHdgs1wtYP3I+Q9zhWaIvEQqHD99wupt75LYbSFVj
Ndm8VnB4Q5VOVqEUHft2ovTAQq5x9phg8w9auMsuzPD4x4Ce5qpWUJ6wCQByvRlwzJCPNGKgWM/Y
wh/cJnI1mXaOizVdP5Ut0quRNL29/uzIgGO+2bqL6KNm8CCBXLU4A0Db12nkCskKfHdv2shl846j
2xl7fxyrA/yifGjCHPcvNO8FPcDTzgHOgxkzuGXndzNE9gkM/6Ir+cH3l4mxOCoVw/P4f7Eqv6Qg
9mS6Gnp6LjVFZt8gLdOpRPsd1oxGXk7Xex5vHMdHexQRkkQ6JJRGwGHXvzXEbE/s1OxBw0soXEOl
kQfyfFGo/I2LzQ94m/1pfXt/oKL5/2XvUCr2zeXATNPqeDjjml6PUaAypMUIjTkreysv+sBLPtOt
VbXsZ7H3+Ney0dZUkVOGymA83I70f5yQpeBKYJuUeV7xWxnIaH1BYpQq3nLQEltCoNxVqRgll1ml
uvLTFBnW7Qy3YuKGwZWFpbNbRC4/SsnjWYuKUEBr6d0BE1clDFzWeB/W3hj+kq9t4h70c0UbGI4C
nUyo97COFDX3hAY5cl59WqRGu8sU0buzFaBoxh7EVkFNi8fxp+fJG7nHwKNJnSZ6KPIMeKifI7gO
qsuIMs/vfNVIMvAL5vEWA2XfzEtpTmztvoH+ow1c0MP1FzTw9GtP/7WMrQaQeakRPOE7EelsNzLJ
h5FYjM+UWLKXXDjUybXPDmwNs2dP4qvBtP4ZhPJwlGhL5z/dkKa+T6f9Lg+Mj/13IMZehyfRB6CO
kg6SUPCTW502t9zBnh5jCXy+qAjn2FKBf6L90e9QsFc+IEsdz70CZiNxjOVuNsxRNXBh2hZY7Mlo
iPYizp/tb2Uq46/zs55K3I74z66s+74ldQ06qKBhgJ3w4XNHnL96mG4z26V24ucRwkBOcZNcXSoi
S6zNWSHJyeznrSVNF6tBBaE1zH6icOpqkIpTr2nRyizmkDRqSPE970n7KpNGcfxNFj6JAb2RtgHJ
FBiZeWS3xqkOwVMVrZdfDlJukl88DxI10dMOYi2BQUlHFCLY+0rCS35tIlXbUib9T6MuDY6vqD2E
bhagX8ylZFmG7zwl6ptP4lHzB9rTC0K/ZFVhr8Pw/eOkUoig0QcfS+GmfJQvZHAGwk5XwW+iB7UQ
3/Z99VW/eKA5RXJOgkA/SPspXueYM78tieKIpdjkw8X60zVqeSg5nB5xsMk8D1OLnn4BeXAd3/Di
mVCVEeO75U5ME3fesQWHIYcx28iLcnA4YoaEJhUtt2T5Z5AnGnwiziEWaEv0J3q2KOvt6zTLvz4h
M//BMWNvgfdyyANeaDXYRGFAUKs5rAxNOSKLMYN012xgLGT3Bf0c9UNT8051uJL0XIXVpPmr4gCf
khtyv5jljbebiPJSUibMsKHADU3zoysktokYhDAZaI8lE2bxmNVd2nssfb7ChDLr+FFeq+F5IiIB
3eJbp/tigTj/Snr6RtyR1ZEZ58yTeoFUt+Gnagdua+m6141nWNeTojxKTS/smm6E+DNKmqS3GlUb
KwCId1MlJ0H7g4gyJndvRpdvJvvQ7ERZF+7+prNSzyWOQ+YVLVLUnPr9s4VeFf4AOBpyPUFoDZIX
/YOVJmY4i8aYHI49rqUhowVFWYXNN5m/1S6V7XfymTCiJPr5Xyscp4+qNmZDKVsqvnnh+cy2TaHL
1RtONyFdrjRsl14lVum0tSM7F2gNddD7sS9qjwJWJdTvwepfFJ5FexJIF42DfkqK/AZie+4n4GtL
xamqR2K1P17PNhC/Gboq6PGXyf9DpunRRfkOXuqBwFzd0tOLCIcSvG4vfehPWU+tPzrpjl/hoAHv
WkQT8+qXm4DdJ+PUgJD43avjgbV2PwffZk3Rnw406UweBoSZgDLtVvPjFL4o7afjquBu+cn4Q9NW
PsF2FPj2SX0bpRi9fahSf8jfsXLwS/1GnRwRDDcwRPjP3M1lhz5aGnSaq/uW719MgKqwqpnS0WaQ
x7bzZjM/Lo6ypvuyq+IWZtO+xwyFbBG0M+IAwyG11DTTNqk48uyxXOhJxhmTNp5oAz8BRshO6YZH
yFGWWlxMKF+1fSC2lrZY3BPou5IrByzYPUk0jGOpbg8kw6wVzfe4zNc6DQEP83789j7eafvqz6pY
Znd0IjdPTvF9R9J+7S0rgrMy8wKtjQDdjqgEUnaSrcBuK0zFpJvwtK2ltaeK42PGa9+x1XecO10L
EdfcainvP6AtLE5Ny9aFeBe8+BZCgGB9SicXtewiedIEFT/k3C2mIuKNTqV0HrhIvKurOl7TudQL
xsKajwAD+RxMbuY51ztPML1/oqoYys6lb0dtKN7jzTQpiv7xzF5R1IYJPqtNjGKWOoahboD542lC
bObZcfWbwCt1eNmfAgXx625G6zprvVN/ggXcu2cr0XkeELbOH8PNnze2Ir44BrYPyP63CLbx1l8s
dwz+ZW+5uOS/EwR/wjWboF5aERfdkgNL/AUnNfmM7C/4W9N519qbMdGtnGxefSperlO4CWASreQ/
lAFMLl64Y6dZB0AoUVjP0ElvYiQwfTeIXBoFSLhBzrK7HUmK5B9DMaMjZ0m7aPZmDJ8v9ZK+iaq+
o/ixXoFh92DRIq+jO5JGmOzUl69HRQirJqKjLLIKVErGoEwOzdsLRoT+oHiMaUv8dtoxEUbJ62ux
pJP1B32/WjNDE4Zx53/Y/ucZj+0QCrrHipLTG1XtQWWrFrzQW9YYL+gowgqRugWGDskGcAP7Wl+S
ySdyNyc7gBOUl5OMIz0rr6N8R8y+OkjDrDB4t/Sv8Ho153EMbLoMuzvf81yoyt6kxMjw7OgP58HK
Xt+yTA3c1oFtnddPGys0qR2kouOfVGDHQNV+A1Fd9OhK7R3uMN3hRdQxKUlzEaD/PngzcWFjDb48
hhX+D6i+8sob8kBgfXE0MIt1DNI2aGlpmZBwJyRsp3DrP+qMycGPLXU5fM2mpbEw8PhgmCmDWfkv
Mpe9hJnIxNJdELnIB1jJKOz8hS5Yap2/zDwspfOAeW0oEsp1vpBhE3yF1Fe0/4ZQKYW00nxW2gww
wFyMOqtgbEe5JbDHh9n+FysxGzMdjlTs6iF68PnrBbkrXbtyugCHpBLZXtySPZPhdVAZjtYWJSFx
fs85tZnn6Pldnc0X9Pd2eL0NLxXfpN7ppzKHPjMWJXkpzFeHHnVkudpM41i5bdlCo5eQH45Uoayt
UOPBZUmoP0m2gNOyW//4hpNLHBoKyqmQanpBpN6hmkS/mEkKCAmyLedf0UFmTJR3+vmQQIUjIh2c
hUTvZubbbIj30vyv2cxbJFd5kRuuWLUZckbWmgOuxdMe3Pz3+t4P7FC25v5JqOkz511GeUtYHwcs
obEByK53C22B3rNo6814Oovj+AvNUlqtCZ29Gq636oPUwZSfhezLKVKN5fWDjLm5B/MD3n8HezhV
Qbk0NZhetbxq3oRgJn/OK5M88ZZ7Iaspg+PFL/lmmUNlpTkYQG33z7bKXlIPrqOQvoJqreE9Vxxu
5txKY5RDeJ6ilwJyDy73B1Ur1C3fKNxMh/Tpk72YAcPcqDs5xniXLNQ0luBaWfplH5wNKdfy5BpX
imJ/WTzvb+0w/SQgz0d0ZhknPUIOqHfBWUwhViceKC/D0oCv+yXv9b5oMHoULBdeA3HceyU1pwde
h2z6e+nFpTuVA/8brRojc5c5jynaKZHYfCxGG6EYqSW4cxfNi0KqmMm5BsGW+mvPfAJwROnN/fJd
iWGKx6pTAi/zHrs0nxckf5KUp3Mlay4R6lyJzal3jDndEIDv2tVVw1qTWwPXx9oVecQkq54DVMkj
mDZy5IEu4K0eqitbyUKWdker6mbf/IrdYI2JL6mq4CAHARaYws65reA/OPERMMYsawRGHaz7yOcl
+t3653MVJ36uXkwvpcFeLyQ7YbdoQ3H90fxrhGHhZons2JZuNmALYKEbzbATh5cqihrK5s2/+seN
cNsJdyudysfeKnlPnpa/OtKA1XA5XQdzOHu0JUyci9L69XBqUfokxFDlbFFB5ny9wP8loMvp7hwy
D9+1IgeDT4Uf93J7gNX57F7dgi55+Zt1nR/uAbdD9VZuUtqHu1OQ/sCxv8+oZ1ZVQcFmJSwJA7FS
UoZU+IrCs7z8QX2j7Gn7JYlslevE38YffDzeh1psBxRzTphliscVaY4uIrn6bgiI+FrjXdUxYZ4K
I8sqTeuS4v9MIYLJMbj8NVfTCuwzJfsrx9NZ5Oj5vvKAlnEc4Jt+VfUyd6i3MDdK5iVJBCB408qf
EbjCw8eRJD5h6Eb5rakK62dZWIXdYhkZ+37fa7gCJsNFKeLm7YLuXro0uc6yv0dBvCK90N5dM5RW
eoHJoQVQsecMVNHpBCou1wVKnWg+dDpLeO170ZwjqHyeHMLw7vPtXA+da4FZ3v4tzlWrwpnmSi0+
KjwVQWXsaX9qZOmXmTnIR7VWbc7mMbcHb2miVOh4vEnY11YaiFGQdibIPtvisPCOsH8xRNNlAwTD
f9m7aVFVdZ4/xcyj5yCqsUtEVXtbdtClfASON5jOESwKQQD7mWfLI6wdPyWXpmVp/QGbuzt6cDa6
YL8/9IHhVBwzQxjbk9U4abUvkLfHFWmsjrT2e0/Q5jJptygOKf4NspdGaQ2kiNU4oDVBnHEqD9Ci
ML3pBKb+XCbfKEeKITTZv0svsR0MkNgtZaHJBQRXEwqS6Cg8ezUbc0WFMJdISD9iyEbdComT3IJ3
sGZYHxunQQsyhwzWEF9ZaumWymQMV71x1jwNXwO2CUYt1rk7zlnk2F6XafT634cTw3FaJBt5Jjxy
7aQdZ3MQqynhXcqXY1J4YlI6JFu/NIQcy9GPiCtDUf4HjPPW9ftE2TpTlof9hBdZ0fprjjwxS9c6
R+DpJn9oRU9QseU00n1c4H6HphdAn6fTBHrO3Nod5oqYTcaRLfJsgetLncpjRFOyxlO3rIkQR1EG
zzRfN78jlhaHmD4kMN2upeoFrPAQHP/wgd5RX6ujrvZmWRT+pb9cVRhsI/bnkMmfoqK2GD+IHWRe
pIHuTKDkkWYdy0r+e8v8+zoHda5z7H7cZYKxlOsLuZlrxqEm41xGBogPaldzKC+wNwYmm43hsQ5y
IYlfiPmAa4GvmBlVCeL0zSSWSd+8quMGPRlMBe6sb0OVf9W4q3nRgpfpdO95NtW0JZHXDyk7UuRl
SB86IBHz+U0qZ5SaQihEXpKbAf2OUGvWgv1+PSx+xZU7nPvVOPhkFYQjFh21YeSDppcquUX+z2By
lgrZutZ/MYmcD7sFV+kSo8QKm614jQW7peoGX5rs6Uck9xPg6ZizXQeuD+3sFNZF42AHzl+3ldkn
GTbrXEV3d8TysoPrv2WhlBn4GiY29ixNc14y9crfr1TrYvrJksyF7/IVZoeU3rAyp25WTJq1j1CB
hGo7NRDflRA8w9Vfgb0UmIo0fIg6W4PS2q7XI4SvV/t3xn3O3qBlCeDsD/afMGdUxDjP77nCkkNJ
C0Vz8VrfG1OD/OCWVXZ833VeWD7iNMP2DAySpfc52UxgyE1Y2Poi6Mk6qIEhS2bGQOv/t00aIqeN
sdsv8tNChdAhQ3oZu2X/x94DqkjAs5N2ejNtBobkPntRoe25+WtpJQWhVVR593shOaAdyTCv+R7N
o4S2k8ru7/JTLZpaYLTba/vXJ5pUFbNmrb4m6Gq1X88KvsesB9xnNfKLlyfmXwjA9NgOzlN242Fg
a3G5tcfzHTw9SkrW2OUFwZEdhKeEqNKO25l76j/oARlqNYQdSE2Zu6VH7fMmBierH+0hGzYWjn0Z
2wCPis9OmCaAr4RmvzzGzXg2+ODDsCXeD1aBl7tav7lArVodJft8oP0b9a2vqsRm2UzIs1bmKdHj
4lJS0RwGtVJ1ZOlzGLt2TN/bOLKc9hzirtryHKQ+/h0o3D3TwFCXydQzrNIae+UhR7A9am3YsCf7
yr4g3qpYolUb3qK6HgK7HyjbCpckGp3ovgem53EIxa3ZyUQFN0FGG6a35Jaiwehm2iSlUgp01LVb
A+H0BQbN3moESMAuf3cti+3MdyANE8CdvkiYGeFSxstkJQS9vtJ4oT2waZibK8gVn2IlIYW5kYxQ
ppSb1ktpiSw/FinplKIkZo/4KjqPoKZdGmKt5K4XhDmWVNMur46QiYg5XSZe+O71v7zVl8xvHTNs
qQYi36u8nyFk2WGWgL6PqGxII6kgiTVScbYHE6a3UI6i7OCgebMeLjbTIWSP/OKYEPlAKwUtSWB0
qaNqk99Hx9ZsDBHBtCm4T7o8sfYRZQZTWyOb0g4vya7rRbsD1tBYzKtWnXFJY0zeCmPQe5bT6/id
MSvlUb+u5Asv3shYH9oQ2Ah3qX+WWCf2kUsS2J/i4lsEmApo+tMvmkxXZYYoCWJoNh6qKXbwaWT3
hkZr/peoVAtFgoktq2pVs53MQOU+vNgsVesP4BRcax+u4jlsmN7ziHGxOXeVlFTPCDi4t8ZDe4G2
YeS1M/Qvx2WrwFe+DBidWLqrVIzCQWUabSngT7S0iyUIb/7nWqrSBvJphGCL/vLoEAsZO3vYvu9b
haFfJEDhtKqJvWlUpZn7h0RRtbA0UbOvTBkxIKIC1dnwXhwYeEkO8tCFwQwkTJ2dGg7CEvFt2Ajv
OmRid7gnN76mpzn94Nmdq0QPRCCYFpsP1jDwTipQvI7MnTKNosgfd28PsmPiVeWKX1Ceqnjj0298
6525+2F92YmRC1eZjFUgvJgtaK52N/q9RyT0Xhe33Q7q0bg7QQENrjnNImCSsNjdQIMFfG8W3i36
pAX4bViQDjCW+z+qO08TxQM2sxK8fVtFR1hbUuLBDoQzALDJqJGCgLDOOHlqbwe7v2pJbnNovlrw
fzJ7+DomwfSm5XEIQTutiRBeXr5k5U/nru1ipgR0G+OWEFSgHyjpVXdeSoDEqnA4qHvT0XUsp+9N
tAE8EM1a/HIQjdkr8fC0yRuTVKbOonqoH6ZyIfhinlHr4DiHPhOTGMPpLPA/nSFkKLdLxMiTex1o
LiaBISYjox7ovvSNzZhCjr7APIUwrb/RNpkfrs4Lpf0GEn6i+vvq1wKVBfhz9GO3SJ8ngCoTvTmn
jWobdVIrQ8FFwfaN3iEPeYDmqRuZhUHFhmX8PBkJxKHdMFIjPXXbVdt0G6IeTwAkkspAT3vtiWLr
+QvqEXXcVHrsA7/huCvuzpl+Jb1avYB7SNXKq0D0PQydcVD/r3DkAkb06x1M1Idw7cm7J8ht8uyl
n1jo033ureY7EEIaXt+q93GCG2g+Lwp1MF9x2By5Pp1amF8i5JL6Zn8lmgP8O4o6gl2nDPKcieuf
lNiHw22RnKxmKFVY9qGj3SaaTo/x0PAv6R1YdW114ud8GNBAt9EU3NsyRevDg7d3u529D2/fbInX
iJGJqGULZRTmwNXfJx9b9TgEbtXxMbsc4BmrzGv6zUC1gI1LchkJjaQ4lMttDrkfxhuAxtyR6vy/
ICdlOxw4kYpV5OVkp/vuG1KRF/6GOoSLdyBDt/hi8Rpm98jvyKbigEVZCCNAC7sJY4A433SWvkAb
pILzso28y+LoR1+1QcZOx/SHnRjV2wnO9oDj4NkXpqdlKm3H2Be2qOTDhw+ql5yfUyGy1L9sBHa0
IKCk87feYV6mlHZJZxCI++SHw5b0fUuvuj9erfySMzgb8MVnJkbmT+gXedYQAk4YFxoM8xHsS3vD
zw2tEC+ck0M4rvD05i5nWr4XGvmq0LIqJXIWntwbpgEPIiMymgzpRGijiLnCRIRo1y1LjxtB+g6D
mh1OleHLpU2t2/JoW2sqo923uhSEdTRaETnpS3E3y61j8DwpfQ9UxCc5mVlgk2qgMquLR6L0DnxE
/Pe47gG4LYssdEMLBtkJQy3R8qZl3M5xkLJqnQzkcoYmlsU1qyZGbrBFnWTGO6p8ypVK36KjULNP
nDjT8wkEKdGr2wT2B3hvdrlxN08XaRlz23QRVDrMkM1jEdqaWQTV48pjpxN33S3fI1hUyl7RdHJe
W914n8t48DeymhEvAgdUlTPRO8/dLvhRTKk8h+dEq6jOnw4H0iFutN4awCF9Pt9bZ9Q1KFIJbSpn
zDql4qyo3o6SDOaEoq65E8Q+s/TDJV82l/GvIp97zkmeB8vA0TrIiuz3rEPcjFY+KqhOUfZHmchC
Eouxqwjo9nbVTo0NwxySrvYTUwpCJzDDJpmZZoTFpGryzQ7Ib0uDq0jyBsDT8mBlAnZsfAx0ZANO
F+rmhjftZYPYt1VL10UUzsQ6nTZucPBeSjBlJnliki8SH/VRvCB4QJb3RlLXn7ytsD7TuzHECMLA
sIOsEmc5HnSoF1hfQg1T7QC5eoqUXZk33QzSGOQF6dumxMRkaCTnpVjbMaDJBfVnoS3eJ6XvLRqb
d2unmmZsRT1wqjJq1E8Mp2TbCPx9JsdRvNjMOlHkgsW4R+ZJQgLCzl09G8c7WckdMvEHhuG5tXKv
NMLWfI4wHksoJMqOCo9UYQfA2mTBkOcSVwwroUquvBprv2Yc40IeK06OW5bZT9ctOyzEJE0NGS/b
HjkY/rgNQjaOadQoAfU3Qb1b3KUk6VSz3xxS2KG8sOdBKMn1eGoNlQDkcXXt88k+fk0HIDm+xZqk
lQBm+hd1fK7odaZCd9k1uj3Sag+KJ6OL6MugeyDNDgFHHTudAEM+led1G3yAQnInNaW290y7WJY6
y1oqCApny8MFBcVteK2F5mBJ6dx6sCnsTdz8oY80ImqQWafmsG/zrjt0VrlXgCTjjf7E00SUbggI
NZykg6aPEPc5ELH+0z5DWvsxdRZsdK2+mGIVKBpsIyqC0U9ee5iNd+R1KmpSTjBqtMevK4TTfF5O
PwVlqLOfslvN3TpZLssz2iP3Dz0H9vZXWRnx67HryolLEpbkWoxvJggg/gRyNiGCw60nUkjKL6uk
Xpcr9HLKYYhKxznnsbyC7HYdlyi3n/IKc+2qC73vD9zi3zE4D65kp4O03cb2oUDp6tfje+PIPnLm
qkjAq4ilhd0VUnI3DX/747rG/bRcFShd2FEvI7RvNSUdvN/msTA7GX79pECiscHbnPez69OgtcDs
CUWw605AkE3g0ebbfSsbOnf9QeNqEoH60vu+rlCcgRy3CXAiVmXNPB93eoiSHlYu7h4qEbtuOUVv
N+OK9nLQbrvIyct4AXpOKOYoz6EArkbyQVQ/i57I0owiScQnY4ancryOim+y1xuHn1x5dsepknRo
EYBm/iNzDPz2FXZ51nHkBTsyvekmEoFiv8y59ccY/CVxxv42zd4EeQdZnGrCeScjRzk3fYFuz3Oo
cC+SMKdqezvPKdCQ8Wvy2ZyigvaOD65qP8INoadnarzCritqTjskEuCLJa6zCmOQXDfeItFBoNgD
1bd53pKgWNG66N2Nxj6N41G1U2YdcXR08jfu4WvNEpWrzhzSOyMDS2zg5xrhbFDcoT8uwkMMDRRv
Sz0JHTH8BhTNO6gPNOvzPDzURc8t1+yAwVOzKDdZhKzrW4wP5JZzTk71l1NTdML/0bfiUV1em83G
oyn1UlImNtDzOV624SKyjlw7YS/26ETW/HGOthw3rIfIwWKIMziX1gDEr44kQ5O6nPue4lidWIpG
4+8GOCgNtSFciJ6g/kP6uzamKExFVJJ/2hA11fC0Yn2DMyJPLVGvDYDrq6Jj6nvatNo0c+hOMzkZ
H5rbsmd2LBqYRMbxFOqCRGzJnuwv5ziOhrMXppMRTjkUSd6eib43cJDD74KO4eFG15YGYZZ2mCrb
QjO6QZuS0YPTh1gavb+8fCP3RsfL2D3q8a4OFouTVuNMf/WRZu9EaV0H26uzMVeaU4v2rgdBTFRm
sRAF7Dza/jkgkHRxMOWqfh0odsoIlZONxO99IGfzp73/XKr+72AZa7qs0l2FBz6z6s4cdLbGo1kY
B24UT8C96xRbCLN8qY+RO4xJdWOCGzwoe4cg81ECsxvZ7yQKI+1QG2AzJTSHGfw8zpPNQA4JC1lz
gwym1HveWPWJOQTq2e1HKHjJgYwjODEhdFDtu9CwGm/sl+i9yntyt/R8GK7GPj8dSboJ8B1zp6Iy
I0ayCncr033IJ91qkyIHuPFPYV9yg8yUk0XG+zpDr+SE3Fink4fWe1eB2s9aOs9LLtXwE47fLM+2
GBfASJOREZzUeGgMEB8S3TozIyDvefQGMR2CH0JCdKLzTu8TlclQzxllrO4zeFmFPflUV8zk2aOa
zWRX1xNLXgEdZ4rAyQZiITTeLwRK7NCME0PHgRD7VI+Gv2vOwVEELN9G6s5AncCYg2N3v2qN25mW
uBezweOLP65QO6BRQGvTJcYFFV3YT3Ag1//lIK3qTlTOSlae1yTZssJB4zAz2+zuCbw58Xq0J0LN
DwPuTKNMl5J0MGEESjAlGUlYEV9Ou94OA67KIWlWFQqUXWuhcqU6azRqxOIAIy1dY+iHVN7Qn6HH
4jfYAfXgL1zLyYmonXuIF8F/2QKORADyVV+8Wu+LS6T5pEVpNLPwElbM8+T3mU0qejD9+uulNa5T
WgvWToQIFhmbDYATZ/KeD97frAmwoycjWa2m5I/aEdLoF4NrTuhQpMzO9/sJTCA44axtsLT28kqs
MMKgleU0IaPnUlSWMxP8Eq7M8kAf6YFFwkdjOlHtPUOVJ2wc+xHlOTz9fxtGcGe4uYyJ9sgXlcvl
j6rhBxemvvU1dC4+5+ResTAkxKYPefcrWEZ5+JsUxByxNaSOUDirKkkAueZn+qXU85KWLScS/wBR
1a7kKFih9bRIsGirRg0/yvE+DPU+xNyLxr/F8qTHxcBkmorC7kjsuHA33aGMyh2FVLN9nBJYuO2S
B15VIXV+sv4e6qJ3fUJpDsUWCikpxP3oi4le3YsjcGArOhiFr6I6P4rjXXTadYsp7lTyqQmfB46U
2nKmRY20d0ZA74zWyPN78lVGMU0sqePyI3a1EhFulwarPewHHXH6v4Z65tU/lqGfwPW3AsxSUthk
j3+wOzj65YYMSnLdMSTeSuf4kdHp7GuLN90YaK2h3G164bJkAjCQsixnYKFlorpsF2HKATKSmDwU
NFpv5DEHEQJxQZqppG2NV21Ok7wMF+x4lXbzgnqzS6G540zmq8vYi8iF+atApZ+lBxS6FsM8gJiP
vf73t8KApnXMad5/Fs0IHahDYi9rOt2cu+1nb5Glg51yekShtuQc87MpmBaUjmNW535KOaeU4Exv
EwTHCQui2i/4sDi0xBZrw3t/eShR115rlMgIkZ+pfnqFJzcAmG7JWCNqBtUX5pyzB92u9iLYi37M
1Y0vtxY/7t1T1zKhsuRBIGBibsI18L+H1k5Qp5Ogu+2+pR8g+h4bcSNOE+V26vdoKpzbyk1wYR0G
yPJNH1C063n4Vq+SzbxfqJFg7EJjtPLa+orxufhVnXzlocO4xTOh5tiJly2lkgpvELKhIRs1cjbQ
+TfpmuTWlaTjW1CcFx9oIwLK3iUjFRzaFOANXOmcWvFMRWQsvfl5eAryHv5fK9GjgNKlyIeGXgNg
FZ9ADSv3VSKTFOYrrrmmNezcyRJIYqn/qd1qA8ou4uykXRhqGP1bdCXmACEEZthezESFzTyu78qI
oFPROQyoEFmf8J1GUivplPQ9wKVmauWe5Mih/9H9Il4C3UrvPKFLhP+WwZr63BxJNixq29FmcSZK
vkmcsQQUvLXzo0S9LEVzf0x3siy5NudwxJNkC3xnmlALQiOaR9Q2VhtSflxLA6i8vzac9zvqT+Dl
0LYPv7P6gI2OfGbrkDigv8YA0YMa/LwGDSTCmiJj9q/MZYUMwwkHEf/Kj7mF/QbiPuCZg097u43o
uDFiz9y9zrkDvMJ553iH7WAqGP1GfvAjIqnt0MqmbiIkGlsaHHZR7YGGlGlA7E41HLhrFLhypV1w
izvZwkdlQMwvtiSnhsEq2sksMool0xVQurtc+f6sR6WZtN2lVXjdGXoDi/Mr2ea3zAPnsOILGe71
qMFefcSDvS1lldN3OqfZGHoYsjQw13Hbhl4t87adse959lGZIfVXQ2s/fuc+QM/Q7KqgR2E9l0Jm
xXsABHvGwA6YPsLyxLV41t9GrOO6ekFKwYs7UqRjoCPl7q0PRE7MJzdBgMJHxBzAyIe8QEfHiTxP
Lkgs9d40UY6aXUpjfrvhV6y6RzwN6yu6kOLVPJJsLFO8wIH3xDhFKS631kvfuskSPG0mz0EQuMf5
KoluJuFZU3JkE7RyLJkDUwK5lZ/9zzbnP291WmCdgrHBad6cYfm9WwVrko5NhjQqhh3NrnDlLFqL
vkJZ+ZoWYT1DZZOmwx4K1gR87L75a9uYBnWfqQJNGnGwZL3HM3vx0VoXkrgNOwh7t5tmqMwQaOcV
/5pwtYCakF5F6Mfrvf0r9ix5L70sXWFctygU0RrGyxgL0tUfHQ/pikkEQ7tAl+rRtaex84VCuxlm
vVfGVQT2KvqIT2F8+TSHuEtdPpMnkaMZnjjZJtkokC/5h94PrKEH/LhgSicWcc4+j8xJPPMMR7yG
UkQLK8F37KpW21CJVzWCWwlCywS4wYUeSQ6cNkklnMoolXTVpA5p4N6qRAxayXA0Dpq/gBQ6t8qp
MjtPt5UXJHT3/d67TjxiDY0wcP13W0qO/aws2HUAE1GThEGSrluDKFsGgKdI2qfpbxrn0PoRN/uy
GjWXZIWaRn43vb4itektzBkQCSG28RIlUSEwy5/I4qbJf0+Il0xoiFvWgHOFN/luRvI42kK7BiGo
I2JznEGM3yl/xTAxHyFqTzajfBgN4z3nWF9qDeu0jFUvMIgHd7YrKN1dTLZcFiERwOg0vBNgx2e8
KtWx0yyahEVsV+NrXuBT3YS8rmDOLcecI9VUHtL3WgK2JcrW1G5Z3h2ho99PbVZ//u+9cw/h+bJV
9Q3JQOm23G+Nhwy720srwOP2+858NvJn+fCDOHoUHPXXbHogTQVJXo5d+VT2mYmB8T8bBh3ZKSlH
3qjwNR9NtM8PUZUDG6IkHgo1gOauIpB/VpeyDzK3WTZvLnToJw1sJ2n79eu9M2csJv8weTM7XFY3
iEs+ujHFlOvRJ6ndNbnQsZdnZX58DeZNrvOOs8uzQwglzKlQTNE5/vsZS0ld69A5xhiVpuow/El8
VYdsGVjF6yKBzbYE3kE1q4WuDWjkKOy1a5uS5ddez1DuSX7pH4+oRTrXAEoeqhJnDfYCn42foGYv
p5DzJaQo3QcK2gmzVPuM/5IoMZwZyR6PVTO/02oB78k7kxHz/jtnS2Ve9lkLp10a7I5CjWsTVq18
QU38gpdOMnpTFWSzbp5z4MxUwBg27IHo3+MnzA9Fjz45+L11BYxQ2OVQ29IlnIVWamTyLnuL5gz5
BzGHDqGN122DRwztHwE4pe5EEvDR+GBSFkp7PB/lnMNUQSDNrz617Lr5wcbnVETt7hOi0uP2FHUL
wht5NjPAtx5eBQwPWm+1UByp+K2ICOoYKgLyjeVb0E7/GQW9GlyA0W1SBeCzpyyyAuPfqSDA+3o5
WaagBLOVCln2YKIpRAcRB4D7o4EC8fQvpuJh7YtHdNeQDF5IlFPl6e/u8sH3A4HMvvs/uIWp4r0Q
H97vU3U69Yc+TxXV1VYLzVVQses+y616Cd5emqyFT9IaBZmQE7b9U5pA1cBiVrp5lORzU70JEy8D
xk3xDbiQILWjvXVt9dYQPvx3PPQdhbtE6YrDp9k+X/G8M+eyBxAXAJUih14CUN4Npn7xq2qYUGCW
8G9/jnd8liHtcXnUvm31TT6ywgsFwNODgmYF+Re0zSrRsuuU9RP28GXVVmN/nMgklIVsFvXXAAZf
JZOpMp7B51efLGapGWj2dcf5su0XU8Sh/LIcpGomzeclbxsddeKzT9OF/kNQneTWD714uDoBTS1P
zdSDCJQjQlbRmp78/OLBRFSVCNmDVy4sKT2k0AmFUcIWFOfiERWKBlio/9rfkzizzeOZ80KtnTJL
GIbKaN11DAkWTUHf5kQksKolaSb3zt5yBamra+aistBsKqVs5hnYXysAoN68FxiWQFREw4+fCtNB
Y4IThvgSm5Y7lRFqZOPXtutyYMMXKjNBcVfmLGhyL3vxbRwYXDVsfnCDFgu8swl4/6pKfeT2I3iM
AtCbBVLR12XifUzAX5oksXk7JBOFy1CQYfPGxfnq9va39exjtCzQujrgAWqHNbWp1exgmcLZZ62s
W1oUIN8YeL0uN+6XnOqc4PXLML3ejho81KIgJbD2aoQv1JtzLDfJ/N1gbUTafghWz+W1LtDfyqaQ
6II59jZb0HN1oYkdAmnHW3NlpQvvp3XQenr8xSQ5RBje/BisRMXyuEsNdZ4+dX+b0dn3ZX7oWCej
jOCN+gjAl5BxxCOYQgXNyukL1nE75MBer8jS/PoRHrV/C1ClYM+0161kOXgOy/a0PqcHUAoyKn89
yAdLwg62VEbu4OkWVZFHXyClYt+F+OZq8lzX8HT9hl4PKzpqnQ1iOn7ksQCS+4Y/UUiUzf7JnM7d
zmFK3y1yocAumWVovI+t/R2it/19NI6swAMcDLIV9IZ4hAyFjRh5I9PLgZQRxC+PVJTSx2uXahp1
n+949oyUi7IJpDHeaczX4o5fKEDYrvP6RiOWKsqg1wTInhuIlysKfMCLXhhuTmvHcSVe56tgj0jp
KfiEXRnZ/I/jPJvXqrtHA96XPTzwI3WvupsYWFZx7b82NmzHPVXxjtIPncqrY3wPrYgvn7X/A10r
GlB6PfpOJWteZ28JqawX82kW8a1GenZ+W+yr1IgWve1qJSdRn6QfkQsL32EEcfu/P9CQw2wWMckx
VlGdu5CSKy0Y7YHVBxx5Tx7KdoHlQwc91Z6KkBdkHAT9/lYpsChqxW0kTBgfDlgvqUkcp+Eb34Ke
VsGzhapoQ4H0TJT7PIC0s3VqGqtQTPf/oa87xUJ2nv7G22BMmQt/oip5FCnO7KfgNVJMFKutlDNa
IdPc4Vvsh0bKUDCvWm84kdfud19nT+OUPfiSOZlBfq2oJpFfGoxBjC4JjGL/ztR4QeugG5L7TsCM
MTGN6U6iZbBiQaRToa1cflHUSvfxUU8WN94KDiPvlBgSiXgtC7YLhWpcB51qHmcWwNagvBFaHSKH
WX2kc3U/yaxYl6oLehRq58CNP2nVkOZt7jJO6KSH/zAJIYoT278Y0tkXj2KeN8PylXw8xaqeRVCm
K1AOT1lsIqkog7kybU5H+4K+PwXD4pFlhmYOs/xJmwzl054y7yfyMIlBH6mOD9/5UkpsFNLwMqUC
wS1GqK9xMZzLCClq6RBv4PIiQBkZNyRLfBtED+wr5UbVkypytxXSLYoE47xvV20pM1ORsQHUmWUN
ZBpSLOBaROl8jyayfNql8LJuUXRmEFGXtirNv/S57vQhhM4571QEkg6xxgwxAsLhXn/tgBZ/tMR6
N0mvbR40RDaKk8J/77jsB9qAqIsS72PsrWHq6V8ee+92VwYAMMx4Jkxqrl26e0Tpr1UW25yiPNFx
6p6gKiWboZ8BNQQm1HhsMKKg942qob22C0FRq6LfGchmRPW9jGP1NbbL3rOVLzWPytmCYh7Be8E5
oWtMbS9hWSn0UgiVeSBvRoLD93Sg56f2SI06arscKaHEkz3k3U/G8E2Uyo1vx9P/uZsjDVWCImak
59kDX2cd8i6gYAiNEr00vY8w5vwN7TYbg6+XK0lFQNeI1ftNWcoqpV993X4HSOMci/XyUvyXJFQO
6HSsh3G921ZUQBAr4rHA1oOCNIzHVewQc4hPd5I8xiJ2UxJPDl73MKt/ACiqeOQK988/NkjKsyz5
OqPYALXrtibbAXfdCVHs87rIXNS8eYRmp6i6D5pqk7w3Qz00PVPSGx3tdYkt5io/VJxho2TUF08M
DPDZ9Z5Sh6+HfJ9WEi0Wbss+EHZdm34tkUi4/HbZnA4bstHbfZu/KaleW6iVlyp7MSd3aCxCOqw4
laJakQ1xo88WD8FnuufyIa5M63DQrQWKQ4CggmCwhTmmj+lEa2YH2HaLHvCaK7OjY2xTz4TyqPhR
iLN891BrD8RjrcT0Y/XaBIWSTbO0HAwvTFZRkRD5bH1id9GVeA3LsQ1zllQaEVwBqTzujnzNts6t
3/aEvzyoZO/HejnbMVatAAHBcYqE2b3OCDPnw68bfb+HCP2lxfCLy1YX/aD5w251Fh1vdS5TBOjp
dMfeyZI2ApzOa2/RDpZRyVjd+A2hK11W9SM/paqMMc8oWitO26vjFB5xnVICetxBDdqPISalMVRu
FAnOzcLRWZ+pYCEoepcPPj1iYCb7MGcKTpot22PRH4qy8Edj4i56r4HfWHezGcSNz4+fyZ+YEnyd
E8M/CRzw0HxOnBZTSW8TnKGqGmzenKzgtvCSfZMb1fxiob3F8/trpgPcvEeWs+A9jaFyJkCnnuEt
H+fA20tm5MFBWGWgaZ4cMvJ76qMj/Pm+XHk2yQa7WaWw+QipTHDizsRDOQmUZXBHx75hfmPeqZPg
83fcyNG2v6O+W1OEqOlqOUd26lr/RUgNvpYexmcmQwInhfy+w/JHyYzv8upXochoDSphgdUJYW/o
J0Fl/gbKyGvqpFqb/O7SjBeRR8loKCoGD5GcHqgVdNGxDn/RFoDIACSMu1wR6jNG8VqXXFkl9Zi+
IuQvF4TwpChoJzC57b/rKauKov/yklQ4drqI21OnW0KDS+9ybLev2OXG/iZ3RaoaC74fzqyt7c9Q
uen+vm/9mthx7OzYYYEE1rfrIqmqE7xinSkgVwuTIETEHD61gkKXg9uRJeQGXMJj0jB+pxtd52WR
z8jHO2eW4/DP/dKs4ac51woZbsjXrtNqcmYmiO2B3jnKtNbdozC7JnKpptxV6aERpgKPZVVAc5Fq
EErWQde2Q8/Hw+d/DynSEJZ4NDY6LQLMRKFpjYdM0KWsH9ink3U1Ta/yZTJlcvjbKsIszrUarTTx
w4mAk9hB8BRQFtk3wLph7aYQO2FCLYuEvN8Urv3QOURHShJBcKSwCV+c1nZufnK+f/IHBzU4ou2X
FWEU3l7I47UIoxOv3Oc8ozopSlidR7BQ3hAfJlaEC2le4RsCtbwrobRdjbCMkG47P3LRgNIHI4Na
qEMY3gDil8di/9j6F8pxwRxEfq0QZdxuzY3tb0t2x5WqVYo84Ron9IIa1/J7+UqcGSPSDtw3RKeY
G4FNeS/K7WY+1hgbG22jifuIbGO9YGclT0WZmkI8ycD0BwRR8mMtkr/o9ixQNN6madBxBrNupRHR
bmD7IfzM+bpuYxFffZjyuRwyPBYQB2S4n5oo5kK/52CpAfaJSv/W0z53kHiqOxLY4nY+7lAGMrD2
wP3EbKrej7HrkAfXKRPrADfZZ9We4GoitMXsw+PYWArqCe+zW5eVijUPE9l+18S9ZX5xu73GwUMu
fOu0EhqRK7EJwVnxnPdnqQsSweex8iYpgrbD4Av9c5ylh6QByPFKVjMMQ1CL5A7CQ/Gw76Fi0BD3
CCDbtOXsl3ww6P1MVh9S2o0FIRx8+I9U7f1mrqwZW7ncAP9I2DhgjvYR6cxwyW4UNJPz00qByr64
eOVzlzJ+h5MS4UjmGlLe7McmBuqAfuc5hcutkYkqeBw6p50vgNMGR5vIllCMaqaSxin/HJbDgsdv
4ET62BrzEn8xwQnrTQ3NMSt/aofIpNkpXTthxsCsQo8b5VcelrfC5nuxchYRUvd9Qa2/hRdg9ddn
dArBL0mvaFJo1+yFWmwj62/iNqBt2ZzQmP6obvIwtm1R68i5ZXtpaqHpgRfc7ER4J/j6AKt0a/Hm
o4iQ7jvrWkcUZb1qa5Ui7l9NNJvRXZaruA/7xpC3+h6qhckWVI1aFPCDFpx6Zrx3Qa0QhwYhNAWZ
yXbnTGKB593x+TJo59Zo2HsTSpfHgozBOE2SCsztr87HuQyNOe4NqOJ1PDAGgwxPmqM83nrW0jDg
a8pUudNFvLmFvBlATbAOqcwwAPDZP5kRxZYHSalDedDwrakY8V4cGZEkFTuGMLKADCZyOEzDth6+
HFwyJIqH8TBD53NsxxuNTM5+jU/n2d7UhsEPzBj+zWJso3XlPwzebtWTMoH/+ix2ZdIrIQxpDNJK
wDwqm83kzz/BbjsTP2dqWaqQXP4ZgDf6LnDrnMJ9DrRqGwud86QbM/VqRLvjb+mc9T41T5XuvHFL
3FfowfvLzxiGXAF8pLi3k7IuftXCuQsXpBFAHbMx2cuFkg7GR4yiFgT8dqC98iVU7qrQ0RLqKLFM
PgGpRBYBlHWpz1LjzMWg4H1c3Iw9brfhgcAvoC/Km5OaM/rIUULWamArQYc2ChOeBYWhdCU/uYVY
1UmILD7t8jADECfsD6hnmyGsgFUo5nQ8WklBMKU1uYnFWynXS2BVFl1gZgfv2bx53jlEkAP2q56X
6RRmrd3+0XEL5nOVTm8x4Km4tW+DjDHqZu9prkZi/06G
`protect end_protected
