-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
suJW/j9guWHUUmKsyS/NeoWc8dsGNoqyyaegf4/drS6TyBXTVNbHNqdgD0iCt3vfOq2TVvT16pyy
PMIkUNwimgKJbquPDOCnZZqf3GrTfQSt5+PdGpLlTAHRiE3oxigQdSeis8z0sRg11/4trrRlcZe2
7wMpG1w8M1xMErc209Y2joP9Xi40RbsYTaOUXm58OQI8lpuuQ2wQr7uP8FAJYPXobjYLGM6wfwQu
V43RjpDKRJEpE4NR4iGWovWZ7mtW1VHlVVxzne2TNn3uQQAYIHacrwFo9wmO+XXraKX6H7CO5dUE
wVDJX8fSHvlCRc/jN1TawJK4/vLztZbK8IPsCg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6160)
`protect data_block
SNk8yulwuNEuISi84yS+5jgqO11pPUKIMfManMROLO4SGtVcI8pBgPMpDP8PGsCDx1fRaPk2LODs
D0LCfWmP+3SWlFlSNASLHT8WGgtJju8Nxxb7qNqFw+HLCxfobXFLb9UMd2K6FnTTuPKXXqin89H8
ajwuz++FQ/syJR4XSfcVHqinFfTqWKvmRjdEHbqRu465UsMfNPqnvM3J+G1+qykCj+vFNI7ndT05
PcuMiFXbLGVFi3yvbVfTNjzu5EzzoWvhsJWWrMB2IjTgLR1n3htMGfgAw7FSF+hpMnECmR1z1IfB
7gxWzdixqBvKjNBr5SAvy6/FMtTtK3/7KvrelKSMizCNFF7byo35fRoZ3LiAbQFtW0AE7RF9fkXn
PbbahAgcL29VCrRd7hcqBQL23wv7+mIAbQfNUcFRMCzoVPT1+LCTHPBop20eN8iI/cT4wIi4N16j
0xsvjlY0dcJj/fecf8d6vxQCvxJ3JU/wOFSZS91sajQLtZbsu4map+hQTMk5O6lAb2BJV31j7Hfc
5qHmuMJXK96X7y7CYlLWlKi6S1WSfULanYWHr9ftZNJSwQBxBQ9ZLBWmtQaV/A/y+QDVPpJwtSmC
hksNm7FkosKxGmliCfwSsxlBAW0OZmXQOazqeWcINeFAtt869JsI8nJKfOvj6mLScClxrl3p/IId
qNr9r/Jd5K70XWSl4Vwbbf1lRZyWS/UUrMkr0wiH6OKg1uTE//n1qb+3hhF+ISptPmhH9rrzh4uf
VQI4lzzZT94vuTJho5WlEFLC9Z4Xl8pU1d+fsSHem5vEsrY3JEhlyCSbID7+r/Rcd9inlIdYVwvh
dM5HDepJ1KMdwT/Md57fsW9f3uZbfAaTmdq7nASl8uuY+8cL7CeGfW7f5fnn5/oXn5f4UYnQT46l
8WzUTd29diuAO2pIPRiywjEokTv6Z+TmYHDr5QNLc7jAPVqPYQnwjVzBXeSjkxDYRjMYdTI3oVeb
OrNN8p6P4Abnso9tfCWv3t4tvDsvguqeLEbpLJR7hwsh9GhmK4MMOf/A7HAaEoo70nX0AfAG2Eo6
HX+vgkO+EpCwCEG7+ceWpv2A4iDBr26iJ/8gmlJ7/v+ftajFQwJwlALVwJ0ZEep3pvZGHRzJNRhm
+I3juMjPFZTxqg/a8/cSPEBwG8zp+/B+oZuaHPrcS8QQ4yXbgqtuI5ZHc3GATAfwpDn53S7eJMA1
lN8GjSrZHvf2Ir3pog01zZM/+X+u/u2kUEP3o/WTCkykNK84IA9mNCL05oON8mRGgSG4xDdEvSDd
nCoSe7CYIBjr4i/lQC8QBdy4q25WwxTXl2C+V5TAPLdPofbKYjcmCWwKv/5WLEdaOBguYVX3UpV0
9IDAM8dX66eM83DkqxTQ+kC1zXRMB7kFcWdYzO7hNMZNaKMPtewk8W1HoaBL9mdKEfNE0wF9K5MH
hc22JOktYHJj4jg7vt7n0iq/QlFWaQENsfoS+IzUQCPLasZjvexDmDMdXSSPZfK3zUlgKLSsUJxP
J43w3pdbGlyQmN7UqlQ/PBFUNxANDKucxsm2fVGQrknalvd6ptebflnmV3lyApnf7AnRGZYP3bTp
6YDIZdGaO9uRTuSz7HpEDh0LOtQRTilr5KT4wo908TPPdz9cYPy6WKMxUPEPNOXXed1oOCGLKfx/
KuZgfEfvYl5XB4Tjbh4Io8pRiXULWwNeFSQ9TqzNa9yX0t1R+F34YrV/GU+2zvzizK9OM1u43Lw4
5dFTYmKxxqKzYOfu7md7MMYj+0m2s2meAX6AddDORBPdEHXFc8rQoDIUE7gLxntyh35/flW/yicl
q/9UYfmNuVBi10AMRTtqTHoz2FeCZVT7OeiKVpnXgcMpmV1krifGu2ebXUk7+u2O9MhVhqnCsvBj
Zj2BXimREgaXxbLjY1lEgnfwcQAsFBFAxViBnK1m/xrwxLTPytPXth00/BRWbMUDVnOMhbC9FQQ7
79GA2Ipg7llN5rg9HeBL7krYqFOAtB0h3WUR6goxdC79hvcnrmEeW9N7/SXArwzuOc0jvbjz5EE0
qdM0CvKtPKwm4ZbQQctkNemFU4cclWr9wD8hoeaK5Py3MR0bcsXK7wRDFYLjJmooasj5AB/ZRvh+
tgh0pjb8l5Ch0xmh5BDbFZ8csl52kuhy2IXL6/EGk9O3Lu9ZtBie3Ho9c7/YLv6UVbOKfLkEmova
pZchUA36JKFhUMivATVNVpBk8/8loiI5DAFynZ7j5GYdKUKp9WYkOh72/FO+aq48+B7MyxJlWco1
E76+Ooh1YRdnkJC54I/KwKFAsAUelbqSfkirzZ37c5WiqABzp8vXoer21YqlypDRrmdQQ+vwEahS
X7VhZO3wGmbcSObDvfVS4csDJLDV835mghXFoGcDe58bvL+Qgrz7FCWfl8mDeoraogt3m0z1usSu
aGwQEw9xKYXr0HOKSd7aIVkBOmHgsT0JAqnoTmcergQgj+xNM3gjBZm+l7OFLwE1pHThcGN8xigv
NA1kU2y91alg+K6Q79hc+UZnyomERf/SiuosepwkD9Odeln2nNqh3GaJsa4Nf87OO3nFK7g6sU+z
Fh6Dgt8UgbmHrvp/h/xL9icuNN43LoOGb+hcbPo54mw0CZ/kwL0bObldTLUXpjctb7h6vnXlouST
nW20B1/6Pzxk9Uq6F+rQEmVFcBdpUtFQha+1pnBwa7m1CgDJKWJgk/Ma3+YcQInZX/cx9KYpn1K3
VkTMQZK9ylYPRo+Pes1X6fjFKqTIDyqmk+fC09YGbM3cCwi2vaDvKT8cHcDgWVC76DXXBqwzMD/5
3oiiFYnqadVB8QmvIgLsv5QwpUAZtTfgBda1Dv/oLDny6UCGOl3IPOjQgPiH8o6nfq1sGEyk0bpi
uzSODvDKg9Dc/QTXexPhCSiEIOWZcYpSL9BD60sFvl1g5jAmWgfkT+x85tud2eCUcygBAE5RIjvB
YheTh0bHufDUH+Rzf3n4dT/D/IbdsG2g0kMkxSthJcIbpYrxynch+gexRzJHH4LHdeWDo5CuRM57
CSCfSTkZZkkD+wBd8s/nl6u1za+mL5ZL9o4AI33eob5SJOmPvbkVBIfMeIpfBJwgEhorlP9SEwWk
a9/SnAOrjR5hgqsHYcb2ZIKoE2jkUECy1Y7GY6BEdzzhaPAW1+oOzTrOjEhpqVbbvV2VPgNwV1uJ
VW5tkQDbESeRcga4Xr3agKQKruqeU7PqW2uhriWWOeWH6SveaIKoLXhv5LeutRQjC6AfMh2dRsyC
RJ3d89fVicG+Yqt1RByB3sEao4vRyFb5A8U1fNOwa1wtQVwzsw77JX7CtnNmfo444BBkH8WqttRV
ySH4lIzUQq4r2jkw8J2wmDBwn/r1nyf8pikxWAlRYTC45cB0+zWpoVsfexQsKahkZGVub17Ui19j
1ltCBK0aGkaooWRO+AeRYPHEDa+bkzrRic4KEYVUuOiMuo+oeeFQs+qjhNP9OmRW/iOBysgi4p9H
e4/zOKMW5M9AcDi4VcRVcR4ZHkgEnPXNi+3gf2NX4dL4cQ7lJrJ8cAsCO790EiLIAfYvVE5SnenX
Q7KuJPW8WBuCf1epxjTyH1w28QrnsFQK0uWXt5LY7UEpZenULF3V5SqejNfN1Pi3OF+2YZcs0Cog
g0bjClOtAzBnBcGXcfoRjyPkZTpnm/x5ehxICUNEP7U/RuCiZQgJoqjJ9px4l4Kziln/4/a/hrNf
wU6u6XoidvLXw1Yknhvn3E/vnhmiTT9cnOXrvOTMm4hEBv5Hx/9Br6qMEHWI/0dQjYcQuRyidrPq
LZ/ZZk01Bt7pr2+l0jqpRtHNWMYQs9TFfFW8iZ+0RzvBi2PDjnw4dATQFr1rLmBj7iArQq8QJ+9n
m8Q1OJeGv3kj4oQTxeatDzZ4pnoee0ZwSR1Tc0VpN5a14pXO6LJJayYqvooXB/i7FFma574GI9bx
GMvHfT8073Ugpt1zaSDfQe/TjcRP5N0wnaD7HeJArfMgjVfWSOZBz9j6nD3IRGNZpGyJfgsVKBPk
mlzlBYBzwFhy82aq0WS5oqAksKyFr14cp9PyHsSgRc1SZ8AX+5L4XfRP/bcloseqhZT1hgl1MNUS
wKd6v3Y90ZyPTw3lEWxUcQgbDcvwOWSfVaXaznYNMkLcTPKnBA6WHn1/HUXfWBIkK4PqfRjz0eUT
WIYX5ddJCrWwOVpLCRQswnguhxLRjZcqdhPR42GxJRSqM4/qv4+PP6NY3leqVW8rrsXOZ2JTsEg8
mqji4PxFFvpJ5hTq4bvjAUqsVqWhLt6BFdNSQgDFRXVktJ+DtQpcxKnoGa+Jc3sfpwP62kLN0dsm
gG0sEzmv3ndWFIFFaaHuGIf3FtHGSjpx7tZkwY3B4x4fC/B8TlI3cjKpn2FP6bnW7bVo7+d7b6xc
9Qc8e+uQ5MwdwiWoLvZieGhfQWna6CHMkQSpKd7NyAphvFuo1ONmGct17p/q8OmEI0knah7bWl4G
VYiFAS5nk7nNkfSsLKUiBY/49XeQEPFwo8tMBoWbKiA0DhB8pWWY6TajNeJzAidiWWyBFEpeEdLO
ulky399qn2/+tmjvewDXeJ5TE9YgckxT4KzcX8SewqZc6ZFkRQgfnTdLFI55nhyyhqKfUhm0E41j
8zpcrSsORKAGm+bnv/OBkd+8JL+RGPqTIkM9hMMSfqPijzauh3v4HZpfZaAlpXf31W6bjKaVWFCr
L10BKMWzWjc8Nri1/gC+O2m3rYZREE/zU5iRaX+Ncf4QD4APXgR3aNaeFdGS/wR+jnB0p81IKeY1
KIn19VW92+zRUJLJlSwy1oCFbMO8kQeeXTbPupYf3YD2pTFMaME0OiOlshKV81zTrau18SpgD/ic
AbguD7YkhWl/7BQiql30GJGbWOhBfxXdIZ/G+mA4p2wrAJIesykVAG33sw21IOjGgQ1YgeWZYLQg
set9K1MOIIexs4Eo7gAaSQ6chXFSRt9m9HIDN5iD31OZ2V6GSBzXhL7uC+H0bEDsEkR0bXVDg652
Jtf6B05vRuO/OBhTR3CpKxUPBW+1/Um/uS6MUzT9wKfdloYv7HndoovZAair2rnqnmA9h+Chj2ic
CwVscBd4ZyizWpf9PRBIJRTzadYLbnbCZCaQpwSf+ywSZyD6IstNUZDLLa0lFG3PI61tPDI8F/xU
PpO7HqyfnWMU6SnvvS+oaLw3zLZMnq46xJKad2Twa46+7efJjX2IL7YCx0AsjDXz5CTxOIFcqPoh
gdTHACoPuB5FoPz2T35aY79l5GrOIAH+NYI+2AOiq2NxoeNiAlMvd8texnVoKTYLnK8114jmn2tE
O4csciX2iknwfbLFaTs3b2baipuwIR0P+/nlJ0lakb7sPnzaDCrqPmG8RKv9FfZDFJQaVQJ/uMXd
OtxTY0lgF780NSAfEJFj6DTYrenA4mxh2ihHQRXHsokg7j4pFA1sy/KCB742VTpjzJ3KnpApDq7z
C8z10Y0aTNX7Hu0RpY1H9EPS2XXdKz0zrXuYtv/ZO0jsNyI5ic7dZUVTAaecN0MHTpC9M5ecLouT
nqXNiTIkict+/y3sgR7mWT0LaQRahVFkPPYHTDj2MwSOqukZW9ahxHqD6maZSO+M0tI/IO+lkzVG
t1N1qa9T4KpwRghwDntWYqnvOK42hvANLW/B0dfRxWf9TFBVuKeyYCke+HHTo3c64EKUy3CdaJl5
k3Ahcfp10BvG2N+wct+LOPuDqBMeCTFg1Q30Nr6FcGbi8ONVG/m3kfXj/6QSRDOQfNjt11w2STUO
Ji9ToQ1o1gF/7WGgV3UV9yStTHrLSuumzDhq8vH51tUyEsW2iAfLaHSSBgjBaKMKM2tI9ibz5gaV
aiizmTyAsj6O1IIivWIErWNSCsdYDs7e4JmJuClUmBjObMh9SLgMl/1dcjTW35StYioy/tdHqIbl
wlk4LLFNhSzyq15saCG4SIsN0W5DzasvL70SxgUiy836i9Bym2k8x7WO2tgS6i9K833L2FeqTbFg
YwS1ykfC0cDtto6McciOttrxAPz1SEl+WvGntou2P4lUebKTxXVKNoc9thDtYlDEyuGww38uiCDZ
hiRW+bdGne+3yOh7fXax/thTcghC/e/a1r4ZLflybyEcYUewfIdDOuOaK0eq7HpnQAN8H4PwPFZz
ca1A4w6KVSk3HUnftA8OLO3o6n/JZeGK1Cqvp4BhsonR8NMOQ4dY2pkiC+HmOpHUm8WWtm84XAvx
MHxAfUXVp7URx9cHR24E5ipEKyjyTnFfJ25wqbY5hxCX01xJgz+8WTfYi0c/XjHZKT0/1j110902
VeZyztXtR82SYnoCYiLlW7HdDGXuupeuG6l8nEaKWEovBXo0mPo1ZmOBBJsoFaTWCje3oIH8tgKz
Fq/iWbWeacpX4psklJ4iRgt1ORtnAD7zhxRwUyS4wP/2p/laaz5ycxNBhXf51TmqzORmvqyjcFDI
0hgGjMPf2NR3FK9BialTez8rAmpjLvx+y1MA5yYwOBw5eAqndQMmKJrBKpyMdJ8qSIxD8AlA2xSO
nu3ZfY9YTEaZ/Q6nlnuONX4dMGCuTAlnfIDGyEfmTyziVJ+eWm760ea7GlZpymMuXTC3g2Pu5UXP
5foImY98d3YSCgj/l2brRthLv+dtq94S+tdgfZreAjfejZqsBYmJ2SdwX1B0MuxzTpkSkYqUtHP2
COyeemT5fEZQd/hANq/S9CUPwK2RcIi9e/vmozjIeVNQqnmXC7rDfu9SgTV6DoRpkFjnGQoVQQPf
4p2qV3V5CDlM+VL0h1t3EF9doJcJOSkwad4fuuUe9yAjnb6MIBzafiDFuuUOK6ulmFzEcNrBTfFp
AHW2+Tf377OcuEPfEPoaxDmNEdFjKBpmGqwtflXDDoAnramfhEzt7gmBB2YWf2dHNy77UF8UrRS5
rx8NifRkpj399r4csfmbNvi5cCBOHLvV8xbiRjq0vKG9gt2kn0tRMgtaZrZwZYvsBybkyfhEmsVY
cBFRNPfmGTRx05cKCKZLjVnpVvR07ElH6wYWdd2nCCzNzCzpm461NsvKIJ/1BXK03UVXknNSqv5c
TxDmbrw5QoVsXvG4lxKQQb5xdABFAe8JtdvVSnGj3NsyKKY/VBY40GARCXZJhD/xG963h4IM3EZ+
UkgGLuPfjNqHo58EnHrvIYlRKjEQc46FDJc1Ms7x2lsoLkJH1EmvSimsNbaT/Cp2gTOKKcSGwnww
HzudOGMRehcEL8h4LzH3Z5uUkR0Y7HvF/lzLstx8DAIHNVZg0pZU2Kg/E1sxY/9mZMOco6ciMqR4
js+g6dlAFqQ+b1sPaLFStSBoptf3u4R0mbPEb+YWSIEy+mGGmj+TdalwRg9DLufVYSThCi7Wray7
LC0SIoPQgyf1SSB/ji6sfwbKlWQiiq4rrm1LsQ6TFMzfalpfA6a45BHEhNNRfgRf5IKOBrWVP4nz
6AZo3IRlog856xE8Oaqxumml7Yqs7IojbrnywbDrTl0ZDk3JSuEIDXT32XK4DMSn1O4WiGZmgHhl
ACzN6jLdqDCo3gWF/kOWVIWjC6SOQEV3ggPcCBFD0lXTBV1wAkDqHotLl860KMOO4TcLhKMwoPng
0gn/WSQ9oVyZq8E6VqBDKj/ulR+4QnuVOsH9alG5VctkMq8ezEGQId3Ud/oDTL9YrNrN0ZpXFmmG
ICpTPxpqjFntkgc45N2yWw0x2r9j+DZOyHCCGfQVPwL0xnTSyos+kXyZVFyCJV00jXH0gCE7Wy4a
ydicP+ELcu45RCBeD9nYN+8fAbfPMzgry3NsgNWTm+KOCVMfcxducatk1K9h3TXqTZoK/BuRb/6D
NDcYiWcqxgzgv0VsxdtDiClWXSQJffNl+JU2Mhafku1ZK/Wvo1HGEvSpl/BzoZ7YN1zE7T1qEwZw
TwErlqvkmrCMP1RiGs9Nc63rtshG8mDeROHLA2Ebb02AnBmjIabEXD0SmO5WtlS9/yZ9EFzURn70
/3bM8wXR452L4VcUl4W79pD56Poq6pAYF1r0HGvqHQBeAkT8yy+WlRWUAbx1VLAJszOOePFDLstg
idH0s80rLvulY8TyE+efjnOhM5ATmF+Ohh+cqcQjEnONI1eIJjuS9pts+1kk4Qf0PA0sPoRv5PmV
Y298eX2FpHwFP+7tTCp4hwkTYU8MlmrQ1Eupq7KN/5KbQg+BlshEd/yuDD1pbvk1olhCViKlrkzn
2tBqgQ==
`protect end_protected
