-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
x8mLXJROchT7YBzK3WrWTyWblJCbgRYpyVkUodA6F9vlg6C875T7IcLp4mTVGt81qqh3nLpTVsOx
6z5gcBucmbEwqCjMOgU3464gAZxZn0G0ES8yuN1lwTpcMgyZjgPFShICY+w1QlylgkkgJ3UebfWK
JPZVZL0zIORmh/I6uGa/yVSRC1ke3kH8X74HPD5AO4ciWeFLzaPDrhcqCrI6qPL+VRgTRp6cV3aj
SQ+jNasuIf26LMLLwRN8iPujMyPLIivUpVjHJNP6VUnjCmY4dn5aiBH3fq1FmB6ztyAqWJAiExbM
WY3P2q8fyydW4WOLLyDGBqaWfRs8RlW2evVeBA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6528)
`protect data_block
vjWP7lRtfWwzxyb83/9uvrnSidZCiARVOXQlIr+46gcW05ILExbBkchBEA5Vy3ysWSA1S5D94sQD
fysifWHPbNxXjXSmXATUc2LTtaceK03n0ovZfmTCZmxLCd/XyeQjieQYarOXCLb2wUR1V6sKISbS
oNr7y020A/A3nuLaAAFp+6T1yP1BXCgy6qXS2KE0zq2lAIrgsRtkw+kWlt5k6wDDxvQdT+xLA4RE
kw52TOL3k5Cb3WAkFWzJ95/B0sLSy8tHJyPi8VUR4UqZuQxhWi6VY0AuZJvZbDAYf4bMsov2VBA1
74RFxD9nhnjMTAGK95GKLFj9F1x9+Kc2HSUa+tfkASEwpdfQCpJLf9367QUBNxKeb6yhXCZ/NKCM
rWfcemsc6EjUSwm2/GoSEXKXGqicWeCBH9m0cNvVT08/1tzVS+khlm7Jm4mPqGVmdtolwDWfrCHu
ILX29nf17llREzi+CR6ihSk+OMoMvaiQ76N8W0T2yi1ZtpkRnNzMob7CmBojpxbk95fzW4Mwc9n2
cACkuDnAQ0Nx08ldrCESp1ixgjE8U/zBYHaaF8BN2mut5iJ9dObSudEMr/YFveXw1vHxky0umHB9
CGgo2CCP6NO/uVzlOi0hy42MYsnJn1KTXNyMjT8mY+dUXxMoLmmMIhB6bPkQJUeKOPmmQZ7Xe4qm
7EC2x4n0k6qJWexNsudWVzipThwgH0fRZKlBS+tIc64CzCq5XtHHp3McLahlqLa5k2ehTZLUKP+v
Wz77c6UA2ZNpQJnNVhpazp+k5ncYtO11kOj+/Wg+gWR4I91tSqk+pMaD7Omshpo5AyVw5h9cq4yO
JG8uSNZ9CYfrbG9Cq6Ba89mqAnm7u8eacMyvCX+9SaELsoeJTu9CCWVtyk6lDVkCGzwJATxXFoVe
2kgWjDPjon4dP51d5PhquzSKfdKMwnEwK1bDrZHfNvtRNFuhA3fY1aCuJ3gTeu1NITkqzGjvXUI8
oSN/i6/KQljdmu06V6Mx5rnwgJffLwtd8+6os5ProDKZuxbtl23flYJrMh9K1WfaOqoHDMaM2Brk
F5nyZUfKMNTjO75xCgmmCwUNnLRLRN3unBgMGOV78F/BW09J+jON7XDYxejaqN4UTsCuv1+ykcbp
Q+ouh1+5WY6LpLF98UsT36l2TZhu99+r4fnF4JHGfvyVQwbZON4KchAwPkaAR+69V+1vVhguC6mS
AGam0MBdPMeiytVbB0GZnAW4P/e1CecqepWzrGFKfzAzkGnSv2OKTYZfFHzC44cza1T+OqIFfzVk
1Gzonuv/DRTKQmxKpaTpeMvptE3qADGW3GnwwPiVaipuaAbQdyWyKRRukHDSlhoPO0YxHT+PvcwO
V9qV2AQCcK+bkru3Yt/acatvrQuprylsrUQCv19K7I2cZk+qzLpKmW5sOOjMi9JbB5sOf+AFHQIk
2eCyv5pH2cKzMpRqqRomTzNA3Lj44yFtSZxA2BYLp1Mudlyftdj/2ApNfZoA/9I6jjeBVUNN6u5U
c0+ueQ+lhbBilIUOAFAn+anfnsBigDpCN5tl1XsC9QuLObYHEnFGQCrws8MTvDjPrn85aAUIVefk
5Y2j7do5PuOFV/JVAAET17aKcH8yae+JYO4lWyybvOubNbvbb/l5c1H46BYegXQVJVuRWxvAXtAw
RnepMRoCeRATtzxyCl3fiqcbL+4HpdTy2zmfpDWhQyzCGkb7a19VAgCy9JofMZNNZDovTMFJ17WG
PjIZ8N9dDhtlMmZSw87io1jgDztgme0hJewUYnDYeONE6s0k28sEZ2DjoOtgFmRIEK4SWZOS+M6e
5An8vJwVADpm9XT5M+J0a3cfP9D1SjpgjeZhF/cWzbLOztbIVKL3y863IGIhdWtmh7axiK29bWw5
XPbM6jVNIP0Eh2aRp8XJfDAV7OgKsAiXy3TmOmMa45upc5fKwYoSoiOKFcoJrecca+aJjh8S2VVZ
Rlgi29/3DMxAM0u/DzSYcywr+GuRpDinmSSk8kYVA6i4WzEhsVx171JELGBzmKfoEVkUv65zGtQd
j8DS1pgSH/G6Pj7UnY37v0ZuczMtx7XzMeSaL4jaPYNzJ4+12GlCd8D1FNejjVNwLyuvhxrxKEXk
t549ameGtz/dp5EGWqIQSjysRZ22YIl0LyQxQu6/qqgZ6IuTXyryGeiWbq7khRhLgIwfPQGNawom
23womZkoUYjOz9I2Hrxx2hU9ELkysF7Wxy86T7t+VuMkCoiu5iKU1LRJZ8JsT5+o4a7gO/ez/n+T
4UEVk8YKkfRHNXs5w42lYhe5GjiecGkPKZa4p3rHOha9v7BflwOftRqzrARD0cJaG9VtsKWKrPVg
gXGQ4SiWAMAU+rFM+8hyHLgMxTl0YfyXb8731B/+KkKRZumBjk0fQAOPbfyGi6nCzvSclW6czP2d
QoKJ2kY6R4sRGU9lsxiW+bfePTDMHSvR82r7vj8MusqpZ/mzMic61Osd6rAyJHng+iitniZBooH4
46uy27GlD/pDOJQ6k5tVa2D46xE7q9m6BsDD8ZgQ+AYDcmG8cfBS3BMzqAQNUo3uVpFr7wu7gFCU
RIgvSES5bXGjgq3vCCvTNisGtvhLPT8b2zZj2gkvGeGtda/DFcpLDKn2OXlgX4X26N6sNXb/gY+Y
mcq3jCCVc2+uhRsnrN4AbDwI683jh7mD2RBmAkFrHsIo+gtz0w7eo5hRNc6cOCB4dML+rrc16eCQ
OrGCNo9JffECfgxvvXhroMbL93SrCIEkCk96j/e8xFEr17j6jLWi2rBzW4QmUBii2X0mdLixPPvv
bf7dKiPJ3uiSADFMWQCNUmzAXu957qveghTqY26E3yhkw4N4gYennav66/KptHB0nPvUwBOECK3a
3TjaX+IaF+1EOzoEAGXTEX280wXqiw5xxn56/cIkb/VILx3xX8asFTjlyFtQoOtFeT0IFuAgO19A
uFANQDv2oyLek430cRAuHP2tizNWVPDmQh6kB0H/RZXZv0mIDR0JUxAq4VO4v7AHpXFdCeaBZuzb
4zKD9n6RRIpThKyGOEPamrq7zfgHibHfrtt1RC5+wgRSNZFok6UDUa5vNjEdIGQ30EQdAxAPkn1m
LZxEaJvHU4WMMQkiR/wz4KWmM+XaGK6QGeATVq679s8KWy64DZaqxdIiHlCa/7spjixyq1aZNdck
DFspVF8NDjE9q4QwKZNgdHqdU5OPu2XAH9NxVoSYZOeYuDJBoeYebHNJrEOk0+Q7gquYxe+4stFI
YIwgW9uL/RMqdw7gtWtIolS2+JiuAUSTiEN8JH1C5+1WofFCbWFxi6GJ8MyNL7PawEcWLnIcNae6
DOZFeZWa6VXjYWwNUxo3o1jMM84bSzkfbA9XoMBpQTY9faGbVT+Q5e645ihcrkkPjIlhUIOhGrge
CuKV1VrWmph8yecI0YbV+heyvw7iayC8HHn5Wb9LKrTWT0M2Al07p2NsW0QbLmGto1avRrNFWWC/
txXrQL31QN9b37eq1DF6OgGxJory8G0Yzl8sf1I6z6/rrmTHmJqAVoo3QyPv02ZVfqwYMYrKPmIo
tEtsRqVs3XnMIiDy5eBOedTX5BwN0LV1d3aKaADz2SU71WldxQhS29zeHegpEDOmt4WC71tj+yX6
dNiI/HXUlAU4N8MjonKQkj33mCoJfBwWAkKTfSmEqapvmPyE876qCoTY/8HGHH2QLH9HFiUSh/gA
wwKzktlzecf80+UwbayIFLTX5r7DHHwkljVfvtXSoMLbRKb/KhWTnPTLu/f1mOkIWHoKmqoOt99T
x9Krd4TJEAuSWgwHdaYsPMAPIX2QbSe5+gtoXY7fFO/VzSq+RZIH1SMrOtd1zd/7bYt1lVzKrACf
/fcEfdZUtMuA67vHU6XC0sdIJIfx5qcM5i+WYpDUKWNUl4E2jw2ZzWah2IiXFY5omAlMlvu48i9P
YDJG3ah88AEKyW5bTHGJburSuLRHEIhfehoFTaN5GFHuLEpGoUWYtosXgl9lTNn4Jj/FhMHgAlJQ
5lJ0a8QrCRLDE9xAazQZg1caPBhf/FzKL3B5xcD7xVbLBP1yH6dCfJWepwpeDPjwLISe6MRwh35m
5NYL1EEBKE5CGL/naK6VWqxgUu0wBxmD8cGa4WLLIuR0zjy0sUGSh5L41SzBSDqQSq/ULgxhtCfp
6ieV9H4dOiav+9G4RVzG+Ahex8XzpoL/yU8wd9jDC2oEQFKTIokElETNNtpdxTV1GoB0f+GlzQi5
IvaaCHyLe14rdWOfCw3OFjBWDn0RYJ7lR95IeoALhjlPLZibJ/JYsCquYEZXmno+OHWSlUQ30U/2
hh7Sb7DhSw4HdsUc/od44TSKGbSsTbMWEbmYqDliSTZH5jHsFgk7sw941scUnp0SSSYbys0AzJ1e
I0bRo6nF2C9KCwKJAA2I0qDypF0wa2SGRXV1JjVegTnGGBhPVdOA7RxptNJZNVXg6+HNO5thv6D1
ZbYyWUIwREPPCKx11RppjD/VPB6PLUZU1lnfTJS/R/eqQqFcihG6fz4UKdD4mgD1NkbuGG1BTiKl
g8gPdSLpKLvi8dRDdPMqDetP9l82lVmnDs+rOMMW03mveQC0VqkWAtwSSm7+qd4ZYlzqPjErDn9I
fZpxz2HqmAAnPssFL3J0nHRn/9fIacl0l7/CfARVJr2OSw0bhvge/CVlwQzyH5sbHGJc7bYOv7qx
cuFtdwWRrw8SitEmz+1czTSrRL+NEjeQUJ9sf6XhjrUrrTRQNxyaEM9eu2fvd5Ukv7R0Opv+7pys
prmQ3+8hUvI3glQ4FZ9Ss2QqEzqIigljMBzhDOwcG/GrexYTAbUuV2VezeBr923tZdw7q9wiB6rT
1FCBPbr16tKKE9IX/9PaG7JlFX9eB9N/Ezsomqw83g0qLSsunQJthaGwPAAFjZ5o0mTg1ZG/FchR
SLvL958czFjFPBZ8mKBCOaVZjx+y2TOF79g+8Pr7TLDBEDN2giRG7yrYAHTi5AcAGgM61WhX8iVg
KlthmQzHiDzbFHF+MiG2WwhsPmQCHrhMTmjZMAU1oTL2jO5KULyQTi8cEmLr8sZRcPRJseV1fxg7
d5EYJMWHj1MLDCRmvIE/sWja44CgCEOwhsSTHeNvMGszXnyfcyIW2xuba3EDw+NDj+gVcRbsZ07M
TwV177zSc1TEJ+ZjJJ5ky/lZgtnodWTfrQB3KMG6+kEPz/k0hBWhlLA7SismXteccWwBZFu3PEDb
F+KpBNS8qOB2NcIg3bACtGhXOKKsnf/dUdNTi2NzSdvK5V6KwaTg3T6nWtqr+KFxaia0ZQWXX7Hz
y0RUpMOxiQgUyahtR7rAui5pxPwe3zAUPVx74yiSzNh2hTR5dHlFD7WaXt8M8vg6zJBn09uiXjrU
jlIFqlhQsdsFWH32PP1sXKbkXdP2yYHrBYN558llRNz35N+/vdUdtFZPGmpOLcruGlJ9NyLRv9hx
cCA6O0BRn6WdmK6x76WY4hquTaFzFxw/XJxx1ExRyzmEo+hN3uFHWoQdrz2pf7MBshR+bv1WoA3L
w225NSMnQ+ANIfXgINvfbE8gJBuqPzOYamtZwez0oC35BgdS7nh3T1aKinEXr9fDwtMeonlmKHV/
Z82tOoO6BrumA5iNEkaYRJYOwpOxUGUQKVIJqFWRXKfOdwrjtmj+7ftlQniTDfNGYTIZlBjAueOq
QE3nXQm3GIXY71+WzCco1uyaSG0HmGHO+hBwlppwOZIuvGeuhHu6Fpp/PtZwdTRHnMrX1V4x8j6M
jmlS1bx1qujFd7FkAkL0Ol0h3pC6ajDaDfWnzgQ/p59rhTNxUFa1kaoMEWYuMqeYICcqPILkEKux
hIlB7/60S/1cF9DjfiLNobAwNcrG4TarGvfm53N0KVcABB5wtxYVrBgrr+4JF+rN2HdWljghVn40
cHXWKBZk+IvGHRg1PcMmZ9g0qBiY668CKivyWYm5xIQz8Kiay6koDWAZu1Lmn2KW1xLW7wteZbzJ
Lrru3SorSa9xQb+af7G/j9wyvVbkPfh8yVoyKIVVn061kJFlsZdM0bxhnOcRb+0hyIpQsjBmEqqV
We2HkygcLiRik4mVamxxFpm6Sl4S7JM5r6uL/7tWJ9LOMLmLG8m9GUmj0AHsrX8sOEiTbAIgqr4y
JitmKnQPgP44bmoliWQ9KaKVDxUK2h+vFr/6dkBtHdOkUDV0FFyIu5MqeJOjkiou5N2ZrLuSH2qX
GJui1/WGQtEJ6kRg0Tl2rkot0NLNQDDIoYHIvd2e57EYvyNRzTXpD+8WdhKEW9chTv1xVS/wJCRs
RERfOMA+peme/JF2KvC1JeoRnkuIpI961Be9892Kq+rvIs0N+p5+tWEVVmkdQU0e2QEUu1iks3bK
iNkX/cusCwFnxqTUODAf1YUWY3miGwNEjBnnRZSKKXsj5MMdryXSCOCssSxYul0SRERpcp+bkoLk
EdvyG9mgloXRnKfWWyQ4aEWfbY8bzJd/G2SDBQCHrACWtOInmfPx9PiGyqEpRZT+YPn2YyNTRJ3m
dGgp61qHhr1X2r4Nsu5HG5hAMFXLxi0HBiUNzYgBSJrgeO77fj/Xs9PUxwnmQQJoVLbdLtlv+32W
lIdYpWgd9q29Vx/oElgq6f4ArVsuD3XiFg4iw5iJJc5qIUfy0hZBfLnMX96QuezgdN1tOh3Jv6Rr
qLXCnINP/mpu7ertui7yIUdnT3vWLv33jH7DLgbYv7pOGCg6cepaGvrQQcWkdO9tsUtnmwroV9nX
73wrW0ZXcptd+fA9+lNeUkTodLAEWFdXC8Oi7+8oN0rnvHAxO0CeE0/2WQK5oswvDiQ7atjjlIAT
m7oA3N2l2exSQ79PuTsCkVeS8z9lnlEpPLMkTdH0belJ7X9r54cGTabIuiHGm1k9TW8jPDJQC9sK
PEBBAWZPPJFeRyQAo74OpDru1p9YI6kl0a84ARvGzKEwXamA6GtzBKanZHck6SYAI4NCnycBO0On
oYn2O2WnN9sk3oMCoTQ5Mvgp+CPDDYjBw9jqYLG80kBsVsmWHD+bLKG4j/cmCUT+qx5SWBxuARYH
NrgNbbmLQCVBQmYiQNEgkMBUmbmStkT1aVAosG0Uq+UVz7LHEsdUhQYFbOzZWutvfYjowQsbWqIS
nhrLXL0UZnP+MprwqImElIVN/nVI2VyCIsMzQGKz4YK7iskK4bPlyQSWRz1iiJOGkccJs5lQMAZs
AzzgDfGMm61Oet6ixaRFNDBPMI3sA8MAXX8aTd6iQPhl5eG9OmWyaHMl0nizD+NTQf5BL5YurMlk
fZtk7QbP4b4gp8XpWOiDkkRdumpWdzX4vaWyjfXwYA4IyEoCcQdRh4lopPC1GPSTCDk5uDKPkOCU
8YhF3DFg+u4BjiNSgQZjDTLF29BCv1O47WqRXsSUtkJ9BRkP0e1bdN/JOrAsrjAjEwuqVwejG8Z8
hUNH0h/jjEEyhbpYLyN4N15o7dshVJRmZthgQrJYVH1WirLbOpxG4T3CK0MfqcL5M8kBLtUHvC+X
HDa3FOjYXsmCIyAii1V36gHwOplrmaGzHVPx8sCoDXE1y2aLpTkxf+RsgA0jll1ikPGtN7yd/HJy
UqoFwhBFKjJ6C50eecGqc3ylHMoGFhwClcnyr46ijH5R+2L8nZUB+Icycb4XXrB+z5yg9URxJzC2
XkW1iUTDXoZVatLwp8afygodDwXyClNAvpFOkw6fntP3jqIEZloDHhK4GgR2y54MHdbl143WF8S7
WcOHKFh2MZoypEU8GxB1IAvmH1tsgpJQqjJPZLIxcw2f3PACqTB20qYz3EkRHPpXQbvFlZUNeB1L
oWFs6ftt+bw0hR1rLvdt8upVjYCNf0tXA/PDtF+1drh1Ao93jSIODoOrjo7Ep6Oi74PNWNGZu3N/
VvRe/OwSNkd4oUeg0M716ra14olgGOwiEdrM+kCECT4qTUGzHXPzDF63P8Woe/M0E15MEuMfk3cU
9H61+aFRrts1LKCnrmJJSNIE1wuxyyQqX07N91y9M5P8Cwv7KpA7mQVcMxgx1UtUnLUcHXQ6v54Y
ifvk4d3y3YgjvbJtfTj5y59kHGSeN8YzLvzCrCXBTho4KIutscUJ1mNZ4YTmo+5k5QJJf9QWjm/c
IOnjFsiL+zsQiwAaiYjYzs/haOl0ecIf414VSOPPAQ+AH+qlODOXXCch2ulfLk0BmpeXDS8nFwii
41nW4iBkusBgkrPLrCnq0BBCziVawWhHcRCSBG3p3+EoTWWsw+FVvXO5tiQ8S/rifPLHTX5+VT0B
/bSZKOZeDUvEf8S4JZREuajGJACTrja+AVggVe8dmd0avqUkvT4j1YNqHG7UXcC1N0QjALO1XJRx
J+iUVT9nm7tkquOlLV0PtP3wlEvphOqzMccw1r55cV/vB/rnJo9HWBgKJrPzQXUARTXU4Cfye02+
6AdUdpjU/G0Q4zVw7dLD6PC8Lctor9RTGiHlyRtuQZh9c+WsDIAe/iFbpTkZePoDqGSs3aZWSHo6
OfV7mEYHlZI9PoviW96FHHi9zGlKimjqpu/wpIqSWozhxeclVTKWw2glhzzfOdCAXzssr+kTVp7p
vODfLrTmnYoqxs80ghE/aUBrCfAfDiLa+8MSC2cflOpgUxkKvIgnRMhoLclILK5tPENgWIa9ZJ/R
Ujxy/TjDyVsVpwANJjfM9vokQz2d74/K7wbMzJYd
`protect end_protected
