��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR���[{�T���CK��TC,���:�
&��d!��]9�'D`�"9 S%�aQ�`!�6������V�W�l�a锦E(�\gC�slu�4U5=1�N�m��l�9ў��P���B�@+yg��=�}|֦���ָJBB����O�� j{(����V� �+X��-�]�0!�G��>�a]��6�,��=0G�L�<�~�|5?����dG5sp��1��c�_�
�Qt�a��F�OG�pZY�c���^;�@ͥ��Y;�k~�S���g��t����W8��E.^�� ҃��W#���tmF�'�~��g�<>%�RN7�l�u'^Z�VHkd�?�	��1>1���s�<}�2AB�|v�7���K����aZyQ��G��L/�m����a��O9lN�|/X/�N�w� ���B�N��v�o�ň�y6�L�B.��n�ա�!�&��D�udK\#��A�_!r4�����74p�t������4?�6y���/�2�����.�=�����
�"-�oO*�nw��a�S,+��\'P��Vc�iL��9�Gf�����ƕ[�]�gі^b�#���t�n|�m��.�S�hx%3�&�Oaÿ�'�M�	�(�,y-�AY�R5+����,C0�b�P62b+۞�ݝ� P�2	�HÄ�;\,&L;�:�������P� L��<�`+���Z!�MWA;��1�w��G����9��w�i��?�Q̈H�
F�dv˥��*3����@4)��|r�mˇ?�1xV�����z4��b��ۍ������=�hFf��˳�-�@M�����e\U6F�G{�S����6��iW��O�Cx�kiY�-{o���7(�i��ϖ'&S���
���5����~�Z�7�tK%4M�*0���e>׺�aG ��>��*,�Oi^1����3OX��l�\�kS&v�g7�ҩ��>9e�-А�(�e-\:�_5�	�M�w�y(@r�7��@�K�w�N;+,�k���ml~I�4���|�+|y�;c~� m�(�680�1����ʮ憁b����5Ky�]~?��R�&��� o��۫�;ֱ"����:�"8�\	�A4ǲ�dw���sZ>�v_�L
��/oW��3/��i矚��3�M\�T�>R��[�m���D���$��j���u?��\%����"�B���{�t)</<��K��C�3��Ĺ�������<���gf:�a��$�B�t�Y<�%OD���53��P^�r�1��� ̍��P��)�����bO�o��nm�.<P3�aR������4��`7�w���#0؆�f�$�&g���r��C��N]�:s~����%z���䍃c�����lm t^n;�9��S��-��1�3��b(gv}�T��V�~*�MĆ����Uь8��\�LO\-����YO [�&��:YD�0�$ۍQQS�9x��a���NwN�g�8�q5��r+�(8}��λ�R����Nf?�Ɓ��1|˧��r�^��p��x�ÿ����B9�. %��(��\�W�$(2�:Ml����@��Y��8=��%�eQ�t��{o1Ö_w8z�ˁ���5�4�ꅠ���̸����[�ǵ��~O&g�b���P��*c�P'�Y�N�5a��a.<�z�%={VD���w7L	���S��Z�1������r'Ҥ��H��7(6^�~��[#K����O�����y�v�0:Pb��H��!�� k,���~,��� ��r�#�&�����Jo��9hI��3o���L{'��U��-:�=,�J�hhl�aڴ��s�./h�8�}�؀�*I�*�)��u�ˮ)���_[��<�#S%��c��W.m���	7akAi������*���|t� ki�m��e��:7p���j�ɥ��+���P_�P�K.H{��@0���E��X�`\m��o�8/��p|G��֙؋���0�4`��z���(�P�԰�k��d�9�Pp���� \�#B��ƕ���A��X�)[��	�zh�i��o����CD��-d;E�j��}�G[���t��[z�qf>)8��y����X�F�;�iT4�S�M���~.���<S��s����EKQ��=t��������"j+�oB-�B���aŽX|�p9Q�t��hoj�z�@�����,�O�f�|if�Z2�朤�te�����Pr=3`C�����)����	�%G;�J�.���d�/�Q,�= �C$�{T� -r�T	�6�M�:�}������w�ѵ��2$�&�4��V�кD\UC[
���wl��^���@�v��{�g/d�=�����>�r�c��gy?<��A�f V�쀙���1~~X�'Qk�c���AjcY2��Zk�/�{_fhg��p"\+��(8�A�nR'�Wx�B����Eve�3)�q��0��<�f["!ű�1�|X+�Z�%��b �yI�b�2�v���mޙ�Gd����@-b�^՛fhd��e�x�W/�Y�=�bo��9�T���ķr>fe�-�e��Nl$�a�)6glfF #[�{j�s+�r(Cn��E+�ڄi�ԅ�K]� �,��5T1j���!jZ�Acu�m&n�/�Zu����y?��'$����P<�	�n�|��si�w�6��'���mw�n!�J���Urꯃ#phQu�`�io�@5}<�&�UY�V$����4�w�r�P�̗-�60Rk �b��Aװ��U��-Z���0�k��k��?GvRc�J$AW��}�'"��F���9D
G'rIV�^vwj�<�	ʧ6��P~)���+��|��l�r�2��Ӹ�.yH��	EOZyu��
<����L�#O&ύ۞�y�T�`T1�E�˛�i#��Â���Z��Tʈna��;	W�J]QU����9�O�m��V���GUw�$Z�C,�q�h;9�+�������� ��,�'��ۈ����6���|L����h��Q��|#%b[ٸ��*�ň�6���a�Y�
�c�����%�佲Ҳ���vX1N�}����e,��D����{&�����d�Z�n����RKQR�F�/2�W5����������gF�0	noa���P�2<�ܠ�8�|�u�
��g{4�<5��;��S﹏\�T���u��+��b%@�k�%sɸ-A^�������Y�7Xk,2�>���;��옖�O�����,��It���_R���gÆ�/E2�`^o��c��5]}����c��=�l����yt}���_�F��7�i�O���)��sσ��%�O���=�C��Meg�(��Js���؉+"�P AK�w�J��@�k���F˲7=�PX�>�4yk@[Nߍ�Q���LsC�tV�� �&�Ӻ�\�~�����Z"��r(���d�L�!�S�ڎt� ��"��J9 �,�"������J<?�f�"��c�tEI-K8�2��JU�6�h�6�a@V_m��H�}�n�/O������0w�"I�*K�E�q�l��C���&ꔄfw��m��)�Ry�Mp�P��nj9�h�K0F�J"]�SG`�xH<����"���lM�s����`e��o.��Z"�j�*>(�����>�6�w�#`N��&�����'��J�*��#���j�����w����.>��G�8��vQy2��!��4."���\|=H�7�q晭>�` ��!�P�涨�� �u�6������Ե��T�g'�2?>��d��h�<D��k����<�D�^�_�gL���:��z*��Kf溇|�vO�1J/%���5���q�m��a3���~@�g�������e�nZ���$���պgjS��#�Cq�M�:ҭM��9����x��J��hVȥ���3��+g�6�����~F;9�"��g^�J���l�=���̶�d;�W�7���X�������Te�R14��̾�8�e�49qY{�t+#O}�!1�9��*T{��i��`�۾�q҂�V�`7wx���w�����ʳ^[�aaP@���eB���[g]������l�|:��5S�>=����%�y<L��9pm�)Jh���r�S������vpq�yKl�4e;�}��]���X���p̑���x�{l�0���?�݄��9��/�7����
u�@�����m��)�O|߼x��)h�� :��������|���Q��4�����6xV�vG�#z�3}Zp�.��*����:���r�5��w��^w~��:���R�I缚��|�Ұ+��)3mǣJg�rG$ߓ�>Y�«��i��i����o(�-O�W��̅1l��:%���-u�+'Z�.�EY��z�7 cS�F,w`���c��e�+�7�|3^���|����;�u�t�2?Hz����@v���,�-�����*�yߠ�|VOI��	i�(�Y6���(U��*>�����x)�ք?U���'M�d���
���:�n���C]Fs��!M�-�R��Ǖ��u�O��c;W����u���,�з�TВ�
J�c{��b`C��=����0�e�&C�q�O5
 �w�{eՍթ}h-,g0}H������-�x�w +DMyg���8�oS��ȵ3�bd:�v�U�f�d��9ێ�@}>J����-i΀r�n�i`^��)�}��%a�֍ro-P��H�P�klր�9i�f-��7���1�>��o��4?#&׫	�e|�[r�ǽ��y}#�k�1R4�!��~Q������h~BK�BOe�R�`w��L�Q����!�y\�{�O�M�a��X	P0�E��� v��'�6hk�
��ϡa�VfQIñ@��W���z%��+4�����\��&�.�-�X��ƺp姴�K���!�Nɬ��:L�_��J�'p��1�k�̽_�Ǧ^f��	@�[�������8�|�Xq��#"�d��9����6�JGj�`�)�T V��g x��p����^\�����lE=�kr\\'���(*���U���-T�_�P�.�w�p��u��J�� t�f��$�͟����"Uֆ;~Rw����F��?x�^�b·IãF�K/ ���Ӧ
�@��2H{�ŴE�0.��>�6Ut��O|�F��I'�CG��>ڝ��{9�#�_@X��#�쫏qs�Y۬t�s'��g��ht}��מ�~Q����%���`���J���a��;![&���yyv�V6����YF���)TV!�˴�im�(��G��9��F�q)dn�CoD6���f�3U��+�+(L/���,86�:��d�}=����0�Ab�[L�����R	�g_�=�"�����*������.c�>�D��m����2�+(@k�ž�D���O �|^�9��7��R��@w��K.�W�_��4,���Ԕ����[��A�I�v$v��ʃI��F�O[��!&�l��1�t3���-x��e�@OB;�!E/C4����ۻ{��+-B[,���loPs~����	���-���aϒhy���Q?�U:�*�Vi[�[��n�9j�����|B��;������^~�և�;K`ݍ�9�5!-��P��rz� �,�L����l��y-�%�jw]�h��4y���y�d�%��:��,Rps!��r�St��ӧ�Pa��wV�je�ػ�S(Q��W{�yH{�%ċ�B�F�U�*���\�x�We/x�b9 �k�)��S�
���9��ب!Mܘ��~r�sU�J��!p�5��R��ެ�0څLk.��,��|s�.���=wY|9%�3����n����3Lr�6+��өH����q��H��AZ��U�`�ZQ�Y�@`�+��MG�Ϧ��v����7���V��p��i��vC'�ۙt��=�p���i����(��uB�4�
o�|VT�,z1?�rߣ8���ǈ9HF
�>�% a�d
o�Ȍ/��8Ϙq����ta��_�M��jqY@u�XV��V�6��jIn��C7����C�&h���A&e=��6�.n����,����ot����=}�k�)-�N$=�J�T�(��\��ta4r���R_V	��ے�;,�-�N��_�F�S���nHCH,oL���TH��U"�k7�^���uX��)_||��#��{����g���x�@ ��J�h���`ȅV}���=u�ރ���T�9����Z
L#|b����5%�B06�J�� ��ZzDN�w�� A�oW=o�%/L��Ƽ��d����zH?ם��>/�Z�]��nڨL�)o�'�k�鷄��Eȥ6��"WQ��}WfX3~Š.��s�b;��ʧRv��2�1r�k��������SA�J��&�1i�m��Uzg�+����G���~��;�R'��Z���L�"@���3�y��ۼ��>˜˞��������Z%�aـ/�<,B�d��x \g�Ƀ�0�uY��\XNe2Tu�DG��!�5x��:��ib<�S�C�:��ؔ$�#W�
�|���z�0����3���̌��?����Cg�px���ΧU�O�η�V��ǎ�h���ĭ����>����h��{�p�ú+��dǂ�
?������Q]�
F�I:��[-���Ġ������
|��H���(+�֓���k]��mCy����%�����bq�m"����]��]��8���H���mm�L_g��fE��/I|��J�!e�'��� p˚�P���9Y�>��N�xܰ�m��OS w��W��5�1a��©��#" 0%��?P�G�b�GMlH�Ժy�~`��!�_>��5�̴E+I��� �)Z�e_�9���]����������Xb�n~�:�ڶ]ܣ��r0-ކ��K�u�>mA��p�k�?�xf�����W�W��q�[�̲0��Ar�O����Ba��&[�'�C\�\�u�roA�g�bR�0/-7�y/�5B���zB������G8��>�Ϗ����2�N:��y�L^Ȅ؝�u��v�m'D�9N6ފ'�ԉ-��oKW,��qr�� D������NfvQء�N�'���	#R�w+5aN���;z�R���K ��p_%0�a_���X�<��a�0UV��B��s�>��®���8��������u�&���dD�X}���D�n�Br���JGB��._q!sn2gT��bb�@r�(C�/��!���X�	��b=~%JN�%��f���/���T��4,`�<���ET�)�ӕ�θs��
������]�Z�
�j��1���B9g�,]�Q�Uk"2�2��+�c�3��pK�2i�������4z���>��e���+�(�k��g��L�up�F�@����4����ztq��>�P�VD�k��#���WI�S��6!��M4�9�����l���5���P��*#j������ʮ�dxjdh��prW�?��2μ7Yp��|k��RC�Μ�&Ub���U�G���];BW˻w���u�U��h��u%3b���yK��b�i�� u�)�q��D�-"�|b�P��0ڃ�U~6�-�Y1����1�6��CHS��Z�����$�I�F�e��Cc߾����`o2�O�-��G�0����P�"���''�B��h������?�"�.� 7��!#�jєo�ZeC��A7�;�|�z�89`
�վ̞��I��:n���y�w@O�yY���G��ck�E3�i��4q�7��0�A��f\|���s��G[�����cv���^��w��]��l�չ0�� Mx��<.$i����Lg��#�2�D�:�~AV1�d*�wp�&��֦o�b��Iw��ƿ���a"A��� �'7��zI�ζ�*M�k��)ӣ�@	$�r��%S	<n�h������zUr�2�v�Ӿ����G�{VVp��7�a�wk��%R.��QǸZ�
r�5�T�ag�j��ʑ����'	~�|��/Ͱ`���-Q�;��.b�86m���8}0~�����T���Q�H���V4���yܴ;>��ݺ �x7@4�5)z\��2�_l��������6�u[���~5\ �S|6��}�%ҫ��w��H�%%�M~D;0����-�b P���+h��Wp,��m?Ѷ�Ǖ��ք�\��@bFp�\n�-�~ �$i�ӱ2���e�?��_o�I��(4tYI���K� ���*@4�C�{br�o�Xk�[�:l{�����g�?y�Vb4b=�	��_��GzPd��}��<( �:a9j4A����%�w9����9�&n�>"��*!�s)���谕i�b�[�o�
^�s��1|۩�*�Y/���颟��ۮ*"����ni�J������#i�
�P}"��g���N!U#���XX�<nq��]�l��Hj i0�W��!���I&��.�
��[ث(F@JN�~ƵME{\�w[h,��q�s��ܠO�UU��x�A�'O���`��&�eէjϋ�a������7��Z����tM��%=�P�!Z�o?}����j=��H[+���D�R�m��긄�-�Y���;��[G/��i#j&wyǡ�޶�L�}��N�׹�T� /�*d�5�������^O�˖�yR���s�;l�6�x��-S����r��a{K��0槒4�=L��`�ri(�!S�߱0��>$�C={�
�3�qi2h`^��F��|4�sP��8D�8k���Iǝ =Z�pC����*�YG�O'��Q/��&�����Ǎ��eG����V;��'�t3��㍛�$`��fGl}=ZE4 ���wş�̻Uu*R�����E�Q�`5pJ�U��
h�r��� �e��]%��Ֆ5�]y�n���5Hy�����Z��|�e>=dj�������ٽn�-