��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR���[{�T���CK��TC,���:�
&��d!��]9�'D`�"9 S%�aQ�`!�6������V�W�l�a锦E(�\gC�slu�4U5=1�N�m��l�9ў��P���B�@+yg+H����Q�����v�Y:���NS�%S��S�@,�^���Y9  ��^�˙��F��3U����`�j0S��O!�,�g�)׃=�`(�h�'{��E~pVʣ�j�)P�J����$4ަ��ܓ�p�V՛���Pu£����![��S�퉞��\�� g�x�> S�
�hN�('�:Z�H9�l��l�#H�>���t���x<��1�^��:�F����~K���糼Tv|�Nos���W�~s	�0~i��LYò.n��BD�;0M1#�]�	�çў�����%R�U�{��bl�j��Wr���[�����v()���MRk���F�Q���Q8}�T�=�[66���ؕ&��։�+��E��;�V<��)k5�t�?}�X��HJ����p�ڝR��SoY�%�֋ϾP��.� �KN�w���d|���L��f]n���8�׬����ň��W�;����7�Y a�ۏ\�m����nx�liA�^Fy�� >���À�x���ռ[���9�ζʔ(�!��Cz��p>�e�G��ѐ�'Ia���~�1�� �1���؝��иG3ao�sv�fǩ�AܬO��SJ���rQL�L ���iA!��k`���#�B�"R��E��wH]f��repRG��,�/ ���'"�ur��k�t�60(�Z�OH�q��ݑ��� ڰ�d�+��D�88_Ϋ>�]�1��<MhO!�b�El4W�a��әN�/���������y?V�a�ܜ�5���xx#˂��a^O,v�kPP�� H��%�ƚټ�m�X�g�
a��u�a��o�Qc(ޚѡv�ڣ�a���d}�ěTwr��m���:�h�>��qB�ٳy�H`�v��I]K�	dȀ�*XX�!=d�6D�qjm9�8�w�+N!ҿG3�C!�Y����x�O�>���,O�a��y��?VOb������2���|�cԇ�J�����K�	f*�@=�,����Z���pG���f6E���1��/8;�TVD�Fc#XS��|��OX�<3Eo{�l�49��x�(YJ统	�t����`ǷEH�D��|�a�00�� Y�Y	��A�`Ҋԑ�@8��
��@L�o����JfW5���n������ʩb�����a4�ɪ��M�`��u�c�7�u��/�L�yD�X����1t�f�i����k�کE9f�i0W!�?��/�	t����庐 b��z`�-��ũ�5C��ڍ��=�h2�$�v�ͭk��N��ΎW�����5k0�_��rbK��-ɯ����OH�5���c>^k���N�>̀���K/_�ݳ���&��=Шm��ƀ�,��Qç�k�J]��X����9c~��d�SpvG�Cr��a�E���(#��y;1���U���S�2�9�Dwd�lC�l`	i�ky{C���,���D�����+��(E��YIcU!��_i�l ��,�~���v&��6�Vi��p��3"��!�Q�;��ʈZ��S��
� ջȋ`J�φ��9eLa�2�B|ܚ(Ѷ�w}� �����ɯ�M� ��������+�ygI����"�d9��sL&����~ 5s��7 �ҹ�{aG*�A�m���6F�����.���d�F�ʁ
�"ߺ�RV��#�-s��y�����[�Е��%Q���S��K�3�
�CY���B�M����#ޠ�m�4��*Ӛ��3���p���b�R'6�*gĭ%�Z�oI��놏�^��Nfc�97Η�w2�:�Z���&F)Q/zo�y��1��/*�֞^Ez�!�vɀ3�bOjպ�'�����{3��P|#!�e~ ѿ�� KI�l�ΐVd���G
^.�M��UEZ�"AD�Џ�"��a�<w��9�׾U`�qV��Z�Յ�-U�&}4�2���X'�-��T�7.K��� o�������%��r� /
����8`��V�ѭg�EjQ[|� �I����NF��U�mr�MDЈ �c�-ࡆX���+��8��7�B���*߸J�K������T< ]�J��e��R�w���L�, a��M�4���	<r����̂U�q^n�?9�/k�2&����!����
m�nF�2-Q�c��m�E�����!/��zg�[X,�R�i��R�/Ivw����u�k�e��}��E��D���]�g���ڧ���-�bD-c�/�<��8�
iyZn��%ٕ����c�|;�gx�A3��Z'r������;Ҿv�ΰ6H�6�p(,�-����)C~�|k7���(U��D(�a�=pG�$�
�S��H~JH'I��y�G�}MzP������F鍧}<�kj1�/dŸ�>����hSc'�sNf����┺8�޴������'y!�G��~�Fh'oEFI����B�vB:�,��8<!H�����3pkN�9v�&�^6��'�I���_�=������yJ�ӒQ�g�I����Ͳڌ
%�Ʈ�>�>����	��� 5�B��:��r1���0����e.�N�2KB������C���̀�s�'z#H����Z�:�/E{+Xyi��Yo\"�y�A�E����@|4v5�jT)��I%^p�ǭ����P�|GYm�rC�'�k`(�Ӈ��#0PIi�lr���o״��S��c�Úς�k�I��k�܂�+;tS���V�