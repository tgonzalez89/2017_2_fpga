-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Ab0RtpaPXNnIYUYbRZ7qsN4jnz5+fCWNoCE1YTgA4E48Ql3FmIqgG369/JoWnAtp5hAdtbKozlB4
jlfCp4NvurN5f0guJMCKdo+whZQ54KzDMf4Eix4o7R9sZJYPcAB4v/QBUjZ7YW8izq+SwRfN4zsp
INpS02ks989eadofWR/3mUdDhs6U/V+f0r+/Zzbn20U4P+Bm7y9IW9yK2+yChoUS688XIteyeK0B
hBe/X8SReMPnvS7Z4D6ja9ljljaIi4g/FTnRADh5WdlVZdPH97WiByRU4w1iSklt+JFecamtneko
InOd/uCJZdWwzv3E1qUukoMhLq/0nucAKkbIUg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 1744)
`protect data_block
8I15cmQOUYXqEZVOWqqnxiVmF1ahSTc89l+ZbaxCRY8wxBF7YwTvXAkgd6t0ZS5tT9TTQLYEEpKn
POKiu3jTfccZtySwnREHIA/Yj0S7KoCY8auRayafAD7Q/VSYfXKSqfsyWpDglwQHdZlH+lXAjg1Q
ONhPQX6hispzi9s+YNTnGtxg8cnDyyGwJ2rIq8481SAiSngCdgABVObYbRU2S/yQGFl9wk3er3EH
6VBO+akbP8Xb9Rus4sOMd8RonlRXF97EAGf6yhTulZdi7DakGikgNaeSs2ieRbkcnz/TvhB4eHU0
no6ET1LWdZgXmeAzllbR2XcUzvGbTFQn26J2ZOKV1Ez/lmPF9CNxaNTtYOtxiF6RzjYw+lY0EShB
KLzuIP1JNGBPbrtwPXS7148wZkbqwGLhxaCoEEBvyLO6H2JhZ/s3EGdhT69UHiAWorGC1z03/nz7
GmOf/KFvHfOCEPhx28x/H1kS+RG6qCTUZHGamq9YuHGCAQykpWtTfFe4TLn4piqNgyIyEThpn9CR
WdznDo3kETjh53vj3P0uVQcyY5VAGMk9DopVdqjVv1ERCWt7mdLYNE5Do+qVwFBv9RJy95pRo0Nt
7MrrZSC8k/LEG1YfPYjfaQExPaVNIBCyGLjCrihOnwRnJibMkLQhD3FX0WZZ1kcKw3Yk4wAkmzkA
H/gQr7jAb8v6qibAxhEps+0Soe1fEoQ5VjKVHFjBA4JMwrVML5yxN6s+62FLJWELhcLhj641blB2
gBlhyX6LmwYC9J1A0jo1oM89p3gmo3RFLp9mfrSfKGwkbKnw79w661NcTr5wptiYbkDNnA1yldX5
r7PKGF1Z6dEkQSwXczIrUEGYbyXu/v/RP5OrmEGGmIJHUI7HNs9ROytngl8kJoTV4n5mTpiBY/2Q
7V3wSULNWqQ//9y8JgRahSmcc6exmH8IL1GX0cy9mch+Wr4W8qxcuocgPeylSnzecyoSRMsDV8tk
t1nISOfOAtCCcsDelXyLDVANRyiwvfr1zce+B6BUrOwkk30G/s5Li2EFl1SKQNoBBAL1d+E9b54G
NrM6dhj2kz6VM08+Fb0Brkg09ab/Vk8TUMjrkTQIGdv2Zqoul95h0WzYg3Y7iQ9RZvNOGKrzPbYC
AXZAAiDjOwf6D+8NUgriMxT8xdkBWp5MzHc2OQnS0P6K2f/qgzJY/MYlyyhLIcCO9F/PQHXAcnHv
6DgMKcB4RbM1Q1eejOsHs52MqWKjspLdowBxI0HEdruPhUC5H5hBgbV1lGZk3RE9d0KCk7zw9K+Z
nAiNoS2FfhP2VHOOFbwBkZAsIg0FkBWh3eQxq7nSpW0+WcxOcxVw16XCvGvq8BBZtH4EU0txqci0
m1Y+0Nja7MPIoRU/PVSMxsraXyUYhZf/BSK1zsKwXEk0wSKLLBX9PizQz5uLyyBrJP/2IHg2UFFo
3tEW6x1rRlDRn/9Sx4erb/U3iygMHsGF0CdJU2Z67MIjMKf66BovnLU2wNsmq+BmTEZXfpOqtWVM
bRHqUtsjvqLa+KIwSb2lCib1NmyI75eFqZShwW3KFV1i40ZTDU0BMHDuE5pn7k23W5tvsM8fFzs9
lP8VpIPvuU39kSETOPh+0QB4kD4P/VMaNeyvepjTc7LzdkWaxSmF1b7hkCI3eRyx9CheEFkpef6I
xUBm7/QxqzC3kyIm90aRdNqZxP/V/HgWH8REh5K8UjWLUDvt+uM+QKB0XrEHKSEzuWW/kDcvY9Nc
Qxcy/QmZjWoufHG020iDhmR6Lxny9vmSONx+PLNCd0GubneJi0RmaW09o8y4Yjzs2lNoPTF+aa6V
1FdkrAAPvknH+aycyTpyweeSX9EcxJt2S/yJo8UV9EKEs9y10u4TvzkS2KBJm4gXft8prJvQEXM3
rIZVrM+6xORfdjyL6JbqkFVi2r2xuXcJMoHdTSVF3V+zbHboH2pvXF1dms/aFm84WZr4YRbIfkPx
kYxqUZfU2VgTqBip5lnAenCwwuMYrQ49z8zoTbAU6e5T+BfD9Zq53EWXxlSWXsMtCoVjB//YJMTd
7M3Hqp5COWVetg/PHob078ef2fbOozUCC2/6LCENnDWOnBicAEa0/EfFAUbOdJpS6LfsqaP0IqYu
IHZsYWGTH/UKxsuI0Y0fg4ciMx7wZ5UUuISJcVrXQcg5wiqXxWQO3q50B+HJONidHeMRIuwIqB7h
/RI+yumrTctiejc1Yst+TEbWNvk5tX8ihf6fCIopcm31lexgqorLAlCv7Yms0I3EEwqTxdFPKSLW
XEz9Ykw3uXY/BB0YGLuhTYqSOEO7BuW419xk/P+oqejLuA==
`protect end_protected
