// Copyright (C) 2017  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Intel and sold by Intel or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// Generated by Quartus Prime Version 16.1.2 Build 203 01/18/2017 SJ Lite Edition
// Created on Tue Jun 20 20:17:09 2017

// synthesis message_off 10175

`timescale 1ns/1ns

module FSM_SPI (
    clock,reset,FIFO_almost_empty,FIFO_empty,Reg_Tx_Empty,
    Reg_Tx_Enable,Mux_Addr_Tx_Sel,Reg_Tx_Req_Data,Reg_Tx_Read_Req);

    input clock;
    input reset;
    input FIFO_almost_empty;
    input FIFO_empty;
    input Reg_Tx_Empty;
    output Reg_Tx_Enable;
    output Mux_Addr_Tx_Sel;
    output Reg_Tx_Req_Data;
    output Reg_Tx_Read_Req;
    reg Reg_Tx_Enable;
    reg Mux_Addr_Tx_Sel;
    reg Reg_Tx_Req_Data;
    reg Reg_Tx_Read_Req;
    reg [3:0] fstate;
    reg [3:0] reg_fstate;
    parameter IDLE=0,A=1,B=2,C=3;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or FIFO_almost_empty or FIFO_empty or Reg_Tx_Empty)
    begin
        if (reset) begin
            reg_fstate <= IDLE;
            Reg_Tx_Enable <= 1'b0;
            Mux_Addr_Tx_Sel <= 1'b0;
            Reg_Tx_Req_Data <= 1'b0;
            Reg_Tx_Read_Req <= 1'b0;
        end
        else begin
            Reg_Tx_Enable <= 1'b0;
            Mux_Addr_Tx_Sel <= 1'b0;
            Reg_Tx_Req_Data <= 1'b0;
            Reg_Tx_Read_Req <= 1'b0;
            case (fstate)
                IDLE: begin
                    if ((FIFO_almost_empty == 1'b0))
                        reg_fstate <= IDLE;
                    else if ((FIFO_almost_empty == 1'b1))
                        reg_fstate <= A;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= IDLE;

                    Mux_Addr_Tx_Sel <= 1'b0;

                    Reg_Tx_Req_Data <= 1'b0;

                    Reg_Tx_Enable <= 1'b0;

                    Reg_Tx_Read_Req <= 1'b0;
                end
                A: begin
                    reg_fstate <= B;

                    Mux_Addr_Tx_Sel <= 1'b0;

                    Reg_Tx_Req_Data <= 1'b0;

                    Reg_Tx_Enable <= 1'b1;

                    Reg_Tx_Read_Req <= 1'b0;
                end
                B: begin
                    if ((Reg_Tx_Empty == 1'b0))
                        reg_fstate <= B;
                    else if ((Reg_Tx_Empty == 1'b1))
                        reg_fstate <= C;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= B;

                    Reg_Tx_Req_Data <= 1'b1;

                    Reg_Tx_Enable <= 1'b0;

                    Reg_Tx_Read_Req <= 1'b0;
                end
                C: begin
                    if ((FIFO_empty == 1'b0))
                        reg_fstate <= B;
                    else if ((FIFO_empty == 1'b1))
                        reg_fstate <= IDLE;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= C;

                    Mux_Addr_Tx_Sel <= 1'b1;

                    Reg_Tx_Req_Data <= 1'b0;

                    Reg_Tx_Enable <= 1'b1;

                    Reg_Tx_Read_Req <= 1'b1;
                end
                default: begin
                    Reg_Tx_Enable <= 1'bx;
                    Mux_Addr_Tx_Sel <= 1'bx;
                    Reg_Tx_Req_Data <= 1'bx;
                    Reg_Tx_Read_Req <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // FSM_gen
